module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \bist_correct[0] ;
 wire \bist_correct[1] ;
 wire \bist_correct[2] ;
 wire \bist_correct[3] ;
 wire \bist_correct[4] ;
 wire \bist_correct[5] ;
 wire \bist_correct[6] ;
 wire \bist_correct[7] ;
 wire \bist_correct_int[0] ;
 wire \bist_correct_int[1] ;
 wire \bist_correct_int[2] ;
 wire \bist_correct_int[3] ;
 wire \bist_correct_int[4] ;
 wire \bist_correct_int[5] ;
 wire \bist_correct_int[6] ;
 wire \bist_correct_int[7] ;
 wire \bist_done[0] ;
 wire \bist_done[1] ;
 wire \bist_done[2] ;
 wire \bist_done[3] ;
 wire \bist_done[4] ;
 wire \bist_done[5] ;
 wire \bist_done[6] ;
 wire \bist_done[7] ;
 wire \bist_done_int[0] ;
 wire \bist_done_int[1] ;
 wire \bist_done_int[2] ;
 wire \bist_done_int[3] ;
 wire \bist_done_int[4] ;
 wire \bist_done_int[5] ;
 wire \bist_done_int[6] ;
 wire \bist_done_int[7] ;
 wire \bist_en[0] ;
 wire \bist_en[1] ;
 wire \bist_en[2] ;
 wire \bist_en[3] ;
 wire \bist_en[4] ;
 wire \bist_en[5] ;
 wire \bist_en[6] ;
 wire \bist_en[7] ;
 wire \bist_en_int[0] ;
 wire \bist_en_int[1] ;
 wire \bist_en_int[2] ;
 wire \bist_en_int[3] ;
 wire \bist_en_int[4] ;
 wire \bist_en_int[5] ;
 wire \bist_en_int[6] ;
 wire \bist_en_int[7] ;
 wire \bist_error[0] ;
 wire \bist_error[1] ;
 wire \bist_error[2] ;
 wire \bist_error[3] ;
 wire \bist_error[4] ;
 wire \bist_error[5] ;
 wire \bist_error[6] ;
 wire \bist_error[7] ;
 wire \bist_error_cnt0[0] ;
 wire \bist_error_cnt0[1] ;
 wire \bist_error_cnt0[2] ;
 wire \bist_error_cnt0[3] ;
 wire \bist_error_cnt0_int[0] ;
 wire \bist_error_cnt0_int[1] ;
 wire \bist_error_cnt0_int[2] ;
 wire \bist_error_cnt0_int[3] ;
 wire \bist_error_cnt1[0] ;
 wire \bist_error_cnt1[1] ;
 wire \bist_error_cnt1[2] ;
 wire \bist_error_cnt1[3] ;
 wire \bist_error_cnt1_int[0] ;
 wire \bist_error_cnt1_int[1] ;
 wire \bist_error_cnt1_int[2] ;
 wire \bist_error_cnt1_int[3] ;
 wire \bist_error_cnt2[0] ;
 wire \bist_error_cnt2[1] ;
 wire \bist_error_cnt2[2] ;
 wire \bist_error_cnt2[3] ;
 wire \bist_error_cnt2_int[0] ;
 wire \bist_error_cnt2_int[1] ;
 wire \bist_error_cnt2_int[2] ;
 wire \bist_error_cnt2_int[3] ;
 wire \bist_error_cnt3[0] ;
 wire \bist_error_cnt3[1] ;
 wire \bist_error_cnt3[2] ;
 wire \bist_error_cnt3[3] ;
 wire \bist_error_cnt3_int[0] ;
 wire \bist_error_cnt3_int[1] ;
 wire \bist_error_cnt3_int[2] ;
 wire \bist_error_cnt3_int[3] ;
 wire \bist_error_cnt4[0] ;
 wire \bist_error_cnt4[1] ;
 wire \bist_error_cnt4[2] ;
 wire \bist_error_cnt4[3] ;
 wire \bist_error_cnt4_int[0] ;
 wire \bist_error_cnt4_int[1] ;
 wire \bist_error_cnt4_int[2] ;
 wire \bist_error_cnt4_int[3] ;
 wire \bist_error_cnt5[0] ;
 wire \bist_error_cnt5[1] ;
 wire \bist_error_cnt5[2] ;
 wire \bist_error_cnt5[3] ;
 wire \bist_error_cnt5_int[0] ;
 wire \bist_error_cnt5_int[1] ;
 wire \bist_error_cnt5_int[2] ;
 wire \bist_error_cnt5_int[3] ;
 wire \bist_error_cnt6[0] ;
 wire \bist_error_cnt6[1] ;
 wire \bist_error_cnt6[2] ;
 wire \bist_error_cnt6[3] ;
 wire \bist_error_cnt6_int[0] ;
 wire \bist_error_cnt6_int[1] ;
 wire \bist_error_cnt6_int[2] ;
 wire \bist_error_cnt6_int[3] ;
 wire \bist_error_cnt7[0] ;
 wire \bist_error_cnt7[1] ;
 wire \bist_error_cnt7[2] ;
 wire \bist_error_cnt7[3] ;
 wire \bist_error_cnt7_int[0] ;
 wire \bist_error_cnt7_int[1] ;
 wire \bist_error_cnt7_int[2] ;
 wire \bist_error_cnt7_int[3] ;
 wire \bist_error_int[0] ;
 wire \bist_error_int[1] ;
 wire \bist_error_int[2] ;
 wire \bist_error_int[3] ;
 wire \bist_error_int[4] ;
 wire \bist_error_int[5] ;
 wire \bist_error_int[6] ;
 wire \bist_error_int[7] ;
 wire \bist_load[0] ;
 wire \bist_load[1] ;
 wire \bist_load[2] ;
 wire \bist_load[3] ;
 wire \bist_load[4] ;
 wire \bist_load[5] ;
 wire \bist_load[6] ;
 wire \bist_load[7] ;
 wire \bist_load_int[0] ;
 wire \bist_load_int[1] ;
 wire \bist_load_int[2] ;
 wire \bist_load_int[3] ;
 wire \bist_load_int[4] ;
 wire \bist_load_int[5] ;
 wire \bist_load_int[6] ;
 wire \bist_load_int[7] ;
 wire bist_rst_n;
 wire \bist_run[0] ;
 wire \bist_run[1] ;
 wire \bist_run[2] ;
 wire \bist_run[3] ;
 wire \bist_run[4] ;
 wire \bist_run[5] ;
 wire \bist_run[6] ;
 wire \bist_run[7] ;
 wire \bist_run_int[0] ;
 wire \bist_run_int[1] ;
 wire \bist_run_int[2] ;
 wire \bist_run_int[3] ;
 wire \bist_run_int[4] ;
 wire \bist_run_int[5] ;
 wire \bist_run_int[6] ;
 wire \bist_run_int[7] ;
 wire \bist_sdi[0] ;
 wire \bist_sdi[1] ;
 wire \bist_sdi[2] ;
 wire \bist_sdi[3] ;
 wire \bist_sdi[4] ;
 wire \bist_sdi[5] ;
 wire \bist_sdi[6] ;
 wire \bist_sdi[7] ;
 wire \bist_sdi_int[0] ;
 wire \bist_sdi_int[1] ;
 wire \bist_sdi_int[2] ;
 wire \bist_sdi_int[3] ;
 wire \bist_sdi_int[4] ;
 wire \bist_sdi_int[5] ;
 wire \bist_sdi_int[6] ;
 wire \bist_sdi_int[7] ;
 wire \bist_sdo[0] ;
 wire \bist_sdo[1] ;
 wire \bist_sdo[2] ;
 wire \bist_sdo[3] ;
 wire \bist_sdo[4] ;
 wire \bist_sdo[5] ;
 wire \bist_sdo[6] ;
 wire \bist_sdo[7] ;
 wire \bist_sdo_int[0] ;
 wire \bist_sdo_int[1] ;
 wire \bist_sdo_int[2] ;
 wire \bist_sdo_int[3] ;
 wire \bist_sdo_int[4] ;
 wire \bist_sdo_int[5] ;
 wire \bist_sdo_int[6] ;
 wire \bist_sdo_int[7] ;
 wire \bist_shift[0] ;
 wire \bist_shift[1] ;
 wire \bist_shift[2] ;
 wire \bist_shift[3] ;
 wire \bist_shift[4] ;
 wire \bist_shift[5] ;
 wire \bist_shift[6] ;
 wire \bist_shift[7] ;
 wire \bist_shift_int[0] ;
 wire \bist_shift_int[1] ;
 wire \bist_shift_int[2] ;
 wire \bist_shift_int[3] ;
 wire \bist_shift_int[4] ;
 wire \bist_shift_int[5] ;
 wire \bist_shift_int[6] ;
 wire \bist_shift_int[7] ;
 wire \cfg_clk_ctrl1[0] ;
 wire \cfg_clk_ctrl1[10] ;
 wire \cfg_clk_ctrl1[11] ;
 wire \cfg_clk_ctrl1[12] ;
 wire \cfg_clk_ctrl1[13] ;
 wire \cfg_clk_ctrl1[14] ;
 wire \cfg_clk_ctrl1[15] ;
 wire \cfg_clk_ctrl1[16] ;
 wire \cfg_clk_ctrl1[17] ;
 wire \cfg_clk_ctrl1[18] ;
 wire \cfg_clk_ctrl1[19] ;
 wire \cfg_clk_ctrl1[1] ;
 wire \cfg_clk_ctrl1[20] ;
 wire \cfg_clk_ctrl1[21] ;
 wire \cfg_clk_ctrl1[22] ;
 wire \cfg_clk_ctrl1[23] ;
 wire \cfg_clk_ctrl1[24] ;
 wire \cfg_clk_ctrl1[25] ;
 wire \cfg_clk_ctrl1[26] ;
 wire \cfg_clk_ctrl1[27] ;
 wire \cfg_clk_ctrl1[28] ;
 wire \cfg_clk_ctrl1[29] ;
 wire \cfg_clk_ctrl1[2] ;
 wire \cfg_clk_ctrl1[30] ;
 wire \cfg_clk_ctrl1[31] ;
 wire \cfg_clk_ctrl1[3] ;
 wire \cfg_clk_ctrl1[4] ;
 wire \cfg_clk_ctrl1[5] ;
 wire \cfg_clk_ctrl1[6] ;
 wire \cfg_clk_ctrl1[7] ;
 wire \cfg_clk_ctrl1[8] ;
 wire \cfg_clk_ctrl1[9] ;
 wire \cfg_clk_ctrl2[0] ;
 wire \cfg_clk_ctrl2[10] ;
 wire \cfg_clk_ctrl2[11] ;
 wire \cfg_clk_ctrl2[12] ;
 wire \cfg_clk_ctrl2[13] ;
 wire \cfg_clk_ctrl2[14] ;
 wire \cfg_clk_ctrl2[15] ;
 wire \cfg_clk_ctrl2[16] ;
 wire \cfg_clk_ctrl2[17] ;
 wire \cfg_clk_ctrl2[18] ;
 wire \cfg_clk_ctrl2[19] ;
 wire \cfg_clk_ctrl2[1] ;
 wire \cfg_clk_ctrl2[20] ;
 wire \cfg_clk_ctrl2[21] ;
 wire \cfg_clk_ctrl2[22] ;
 wire \cfg_clk_ctrl2[23] ;
 wire \cfg_clk_ctrl2[24] ;
 wire \cfg_clk_ctrl2[25] ;
 wire \cfg_clk_ctrl2[26] ;
 wire \cfg_clk_ctrl2[27] ;
 wire \cfg_clk_ctrl2[28] ;
 wire \cfg_clk_ctrl2[29] ;
 wire \cfg_clk_ctrl2[2] ;
 wire \cfg_clk_ctrl2[30] ;
 wire \cfg_clk_ctrl2[31] ;
 wire \cfg_clk_ctrl2[3] ;
 wire \cfg_clk_ctrl2[4] ;
 wire \cfg_clk_ctrl2[5] ;
 wire \cfg_clk_ctrl2[6] ;
 wire \cfg_clk_ctrl2[7] ;
 wire \cfg_clk_ctrl2[8] ;
 wire \cfg_clk_ctrl2[9] ;
 wire lbist_clk;
 wire \mem1_addr_a[10] ;
 wire \mem1_addr_a[2] ;
 wire \mem1_addr_a[3] ;
 wire \mem1_addr_a[4] ;
 wire \mem1_addr_a[5] ;
 wire \mem1_addr_a[6] ;
 wire \mem1_addr_a[7] ;
 wire \mem1_addr_a[8] ;
 wire \mem1_addr_a[9] ;
 wire \mem1_addr_b[10] ;
 wire \mem1_addr_b[2] ;
 wire \mem1_addr_b[3] ;
 wire \mem1_addr_b[4] ;
 wire \mem1_addr_b[5] ;
 wire \mem1_addr_b[6] ;
 wire \mem1_addr_b[7] ;
 wire \mem1_addr_b[8] ;
 wire \mem1_addr_b[9] ;
 wire mem1_cen_a;
 wire mem1_cen_b;
 wire mem1_clk_a;
 wire mem1_clk_b;
 wire \mem1_din_b[0] ;
 wire \mem1_din_b[10] ;
 wire \mem1_din_b[11] ;
 wire \mem1_din_b[12] ;
 wire \mem1_din_b[13] ;
 wire \mem1_din_b[14] ;
 wire \mem1_din_b[15] ;
 wire \mem1_din_b[16] ;
 wire \mem1_din_b[17] ;
 wire \mem1_din_b[18] ;
 wire \mem1_din_b[19] ;
 wire \mem1_din_b[1] ;
 wire \mem1_din_b[20] ;
 wire \mem1_din_b[21] ;
 wire \mem1_din_b[22] ;
 wire \mem1_din_b[23] ;
 wire \mem1_din_b[24] ;
 wire \mem1_din_b[25] ;
 wire \mem1_din_b[26] ;
 wire \mem1_din_b[27] ;
 wire \mem1_din_b[28] ;
 wire \mem1_din_b[29] ;
 wire \mem1_din_b[2] ;
 wire \mem1_din_b[30] ;
 wire \mem1_din_b[31] ;
 wire \mem1_din_b[3] ;
 wire \mem1_din_b[4] ;
 wire \mem1_din_b[5] ;
 wire \mem1_din_b[6] ;
 wire \mem1_din_b[7] ;
 wire \mem1_din_b[8] ;
 wire \mem1_din_b[9] ;
 wire \mem1_dout_a[0] ;
 wire \mem1_dout_a[10] ;
 wire \mem1_dout_a[11] ;
 wire \mem1_dout_a[12] ;
 wire \mem1_dout_a[13] ;
 wire \mem1_dout_a[14] ;
 wire \mem1_dout_a[15] ;
 wire \mem1_dout_a[16] ;
 wire \mem1_dout_a[17] ;
 wire \mem1_dout_a[18] ;
 wire \mem1_dout_a[19] ;
 wire \mem1_dout_a[1] ;
 wire \mem1_dout_a[20] ;
 wire \mem1_dout_a[21] ;
 wire \mem1_dout_a[22] ;
 wire \mem1_dout_a[23] ;
 wire \mem1_dout_a[24] ;
 wire \mem1_dout_a[25] ;
 wire \mem1_dout_a[26] ;
 wire \mem1_dout_a[27] ;
 wire \mem1_dout_a[28] ;
 wire \mem1_dout_a[29] ;
 wire \mem1_dout_a[2] ;
 wire \mem1_dout_a[30] ;
 wire \mem1_dout_a[31] ;
 wire \mem1_dout_a[3] ;
 wire \mem1_dout_a[4] ;
 wire \mem1_dout_a[5] ;
 wire \mem1_dout_a[6] ;
 wire \mem1_dout_a[7] ;
 wire \mem1_dout_a[8] ;
 wire \mem1_dout_a[9] ;
 wire \mem1_mask_b[0] ;
 wire \mem1_mask_b[1] ;
 wire \mem1_mask_b[2] ;
 wire \mem1_mask_b[3] ;
 wire mem1_web_b;
 wire \mem2_addr_a[10] ;
 wire \mem2_addr_a[2] ;
 wire \mem2_addr_a[3] ;
 wire \mem2_addr_a[4] ;
 wire \mem2_addr_a[5] ;
 wire \mem2_addr_a[6] ;
 wire \mem2_addr_a[7] ;
 wire \mem2_addr_a[8] ;
 wire \mem2_addr_a[9] ;
 wire \mem2_addr_b[10] ;
 wire \mem2_addr_b[2] ;
 wire \mem2_addr_b[3] ;
 wire \mem2_addr_b[4] ;
 wire \mem2_addr_b[5] ;
 wire \mem2_addr_b[6] ;
 wire \mem2_addr_b[7] ;
 wire \mem2_addr_b[8] ;
 wire \mem2_addr_b[9] ;
 wire mem2_cen_a;
 wire mem2_cen_b;
 wire mem2_clk_a;
 wire mem2_clk_b;
 wire \mem2_din_b[0] ;
 wire \mem2_din_b[10] ;
 wire \mem2_din_b[11] ;
 wire \mem2_din_b[12] ;
 wire \mem2_din_b[13] ;
 wire \mem2_din_b[14] ;
 wire \mem2_din_b[15] ;
 wire \mem2_din_b[16] ;
 wire \mem2_din_b[17] ;
 wire \mem2_din_b[18] ;
 wire \mem2_din_b[19] ;
 wire \mem2_din_b[1] ;
 wire \mem2_din_b[20] ;
 wire \mem2_din_b[21] ;
 wire \mem2_din_b[22] ;
 wire \mem2_din_b[23] ;
 wire \mem2_din_b[24] ;
 wire \mem2_din_b[25] ;
 wire \mem2_din_b[26] ;
 wire \mem2_din_b[27] ;
 wire \mem2_din_b[28] ;
 wire \mem2_din_b[29] ;
 wire \mem2_din_b[2] ;
 wire \mem2_din_b[30] ;
 wire \mem2_din_b[31] ;
 wire \mem2_din_b[3] ;
 wire \mem2_din_b[4] ;
 wire \mem2_din_b[5] ;
 wire \mem2_din_b[6] ;
 wire \mem2_din_b[7] ;
 wire \mem2_din_b[8] ;
 wire \mem2_din_b[9] ;
 wire \mem2_dout_a[0] ;
 wire \mem2_dout_a[10] ;
 wire \mem2_dout_a[11] ;
 wire \mem2_dout_a[12] ;
 wire \mem2_dout_a[13] ;
 wire \mem2_dout_a[14] ;
 wire \mem2_dout_a[15] ;
 wire \mem2_dout_a[16] ;
 wire \mem2_dout_a[17] ;
 wire \mem2_dout_a[18] ;
 wire \mem2_dout_a[19] ;
 wire \mem2_dout_a[1] ;
 wire \mem2_dout_a[20] ;
 wire \mem2_dout_a[21] ;
 wire \mem2_dout_a[22] ;
 wire \mem2_dout_a[23] ;
 wire \mem2_dout_a[24] ;
 wire \mem2_dout_a[25] ;
 wire \mem2_dout_a[26] ;
 wire \mem2_dout_a[27] ;
 wire \mem2_dout_a[28] ;
 wire \mem2_dout_a[29] ;
 wire \mem2_dout_a[2] ;
 wire \mem2_dout_a[30] ;
 wire \mem2_dout_a[31] ;
 wire \mem2_dout_a[3] ;
 wire \mem2_dout_a[4] ;
 wire \mem2_dout_a[5] ;
 wire \mem2_dout_a[6] ;
 wire \mem2_dout_a[7] ;
 wire \mem2_dout_a[8] ;
 wire \mem2_dout_a[9] ;
 wire \mem2_mask_b[0] ;
 wire \mem2_mask_b[1] ;
 wire \mem2_mask_b[2] ;
 wire \mem2_mask_b[3] ;
 wire mem2_web_b;
 wire \mem3_addr_a[10] ;
 wire \mem3_addr_a[2] ;
 wire \mem3_addr_a[3] ;
 wire \mem3_addr_a[4] ;
 wire \mem3_addr_a[5] ;
 wire \mem3_addr_a[6] ;
 wire \mem3_addr_a[7] ;
 wire \mem3_addr_a[8] ;
 wire \mem3_addr_a[9] ;
 wire \mem3_addr_b[10] ;
 wire \mem3_addr_b[2] ;
 wire \mem3_addr_b[3] ;
 wire \mem3_addr_b[4] ;
 wire \mem3_addr_b[5] ;
 wire \mem3_addr_b[6] ;
 wire \mem3_addr_b[7] ;
 wire \mem3_addr_b[8] ;
 wire \mem3_addr_b[9] ;
 wire mem3_cen_a;
 wire mem3_cen_b;
 wire mem3_clk_a;
 wire mem3_clk_b;
 wire \mem3_din_b[0] ;
 wire \mem3_din_b[10] ;
 wire \mem3_din_b[11] ;
 wire \mem3_din_b[12] ;
 wire \mem3_din_b[13] ;
 wire \mem3_din_b[14] ;
 wire \mem3_din_b[15] ;
 wire \mem3_din_b[16] ;
 wire \mem3_din_b[17] ;
 wire \mem3_din_b[18] ;
 wire \mem3_din_b[19] ;
 wire \mem3_din_b[1] ;
 wire \mem3_din_b[20] ;
 wire \mem3_din_b[21] ;
 wire \mem3_din_b[22] ;
 wire \mem3_din_b[23] ;
 wire \mem3_din_b[24] ;
 wire \mem3_din_b[25] ;
 wire \mem3_din_b[26] ;
 wire \mem3_din_b[27] ;
 wire \mem3_din_b[28] ;
 wire \mem3_din_b[29] ;
 wire \mem3_din_b[2] ;
 wire \mem3_din_b[30] ;
 wire \mem3_din_b[31] ;
 wire \mem3_din_b[3] ;
 wire \mem3_din_b[4] ;
 wire \mem3_din_b[5] ;
 wire \mem3_din_b[6] ;
 wire \mem3_din_b[7] ;
 wire \mem3_din_b[8] ;
 wire \mem3_din_b[9] ;
 wire \mem3_dout_a[0] ;
 wire \mem3_dout_a[10] ;
 wire \mem3_dout_a[11] ;
 wire \mem3_dout_a[12] ;
 wire \mem3_dout_a[13] ;
 wire \mem3_dout_a[14] ;
 wire \mem3_dout_a[15] ;
 wire \mem3_dout_a[16] ;
 wire \mem3_dout_a[17] ;
 wire \mem3_dout_a[18] ;
 wire \mem3_dout_a[19] ;
 wire \mem3_dout_a[1] ;
 wire \mem3_dout_a[20] ;
 wire \mem3_dout_a[21] ;
 wire \mem3_dout_a[22] ;
 wire \mem3_dout_a[23] ;
 wire \mem3_dout_a[24] ;
 wire \mem3_dout_a[25] ;
 wire \mem3_dout_a[26] ;
 wire \mem3_dout_a[27] ;
 wire \mem3_dout_a[28] ;
 wire \mem3_dout_a[29] ;
 wire \mem3_dout_a[2] ;
 wire \mem3_dout_a[30] ;
 wire \mem3_dout_a[31] ;
 wire \mem3_dout_a[3] ;
 wire \mem3_dout_a[4] ;
 wire \mem3_dout_a[5] ;
 wire \mem3_dout_a[6] ;
 wire \mem3_dout_a[7] ;
 wire \mem3_dout_a[8] ;
 wire \mem3_dout_a[9] ;
 wire \mem3_mask_b[0] ;
 wire \mem3_mask_b[1] ;
 wire \mem3_mask_b[2] ;
 wire \mem3_mask_b[3] ;
 wire mem3_web_b;
 wire \mem4_addr_a[10] ;
 wire \mem4_addr_a[2] ;
 wire \mem4_addr_a[3] ;
 wire \mem4_addr_a[4] ;
 wire \mem4_addr_a[5] ;
 wire \mem4_addr_a[6] ;
 wire \mem4_addr_a[7] ;
 wire \mem4_addr_a[8] ;
 wire \mem4_addr_a[9] ;
 wire \mem4_addr_b[10] ;
 wire \mem4_addr_b[2] ;
 wire \mem4_addr_b[3] ;
 wire \mem4_addr_b[4] ;
 wire \mem4_addr_b[5] ;
 wire \mem4_addr_b[6] ;
 wire \mem4_addr_b[7] ;
 wire \mem4_addr_b[8] ;
 wire \mem4_addr_b[9] ;
 wire mem4_cen_a;
 wire mem4_cen_b;
 wire mem4_clk_a;
 wire mem4_clk_b;
 wire \mem4_din_b[0] ;
 wire \mem4_din_b[10] ;
 wire \mem4_din_b[11] ;
 wire \mem4_din_b[12] ;
 wire \mem4_din_b[13] ;
 wire \mem4_din_b[14] ;
 wire \mem4_din_b[15] ;
 wire \mem4_din_b[16] ;
 wire \mem4_din_b[17] ;
 wire \mem4_din_b[18] ;
 wire \mem4_din_b[19] ;
 wire \mem4_din_b[1] ;
 wire \mem4_din_b[20] ;
 wire \mem4_din_b[21] ;
 wire \mem4_din_b[22] ;
 wire \mem4_din_b[23] ;
 wire \mem4_din_b[24] ;
 wire \mem4_din_b[25] ;
 wire \mem4_din_b[26] ;
 wire \mem4_din_b[27] ;
 wire \mem4_din_b[28] ;
 wire \mem4_din_b[29] ;
 wire \mem4_din_b[2] ;
 wire \mem4_din_b[30] ;
 wire \mem4_din_b[31] ;
 wire \mem4_din_b[3] ;
 wire \mem4_din_b[4] ;
 wire \mem4_din_b[5] ;
 wire \mem4_din_b[6] ;
 wire \mem4_din_b[7] ;
 wire \mem4_din_b[8] ;
 wire \mem4_din_b[9] ;
 wire \mem4_dout_a[0] ;
 wire \mem4_dout_a[10] ;
 wire \mem4_dout_a[11] ;
 wire \mem4_dout_a[12] ;
 wire \mem4_dout_a[13] ;
 wire \mem4_dout_a[14] ;
 wire \mem4_dout_a[15] ;
 wire \mem4_dout_a[16] ;
 wire \mem4_dout_a[17] ;
 wire \mem4_dout_a[18] ;
 wire \mem4_dout_a[19] ;
 wire \mem4_dout_a[1] ;
 wire \mem4_dout_a[20] ;
 wire \mem4_dout_a[21] ;
 wire \mem4_dout_a[22] ;
 wire \mem4_dout_a[23] ;
 wire \mem4_dout_a[24] ;
 wire \mem4_dout_a[25] ;
 wire \mem4_dout_a[26] ;
 wire \mem4_dout_a[27] ;
 wire \mem4_dout_a[28] ;
 wire \mem4_dout_a[29] ;
 wire \mem4_dout_a[2] ;
 wire \mem4_dout_a[30] ;
 wire \mem4_dout_a[31] ;
 wire \mem4_dout_a[3] ;
 wire \mem4_dout_a[4] ;
 wire \mem4_dout_a[5] ;
 wire \mem4_dout_a[6] ;
 wire \mem4_dout_a[7] ;
 wire \mem4_dout_a[8] ;
 wire \mem4_dout_a[9] ;
 wire \mem4_mask_b[0] ;
 wire \mem4_mask_b[1] ;
 wire \mem4_mask_b[2] ;
 wire \mem4_mask_b[3] ;
 wire mem4_web_b;
 wire \mem5_addr_a[2] ;
 wire \mem5_addr_a[3] ;
 wire \mem5_addr_a[4] ;
 wire \mem5_addr_a[5] ;
 wire \mem5_addr_a[6] ;
 wire \mem5_addr_a[7] ;
 wire \mem5_addr_a[8] ;
 wire \mem5_addr_a[9] ;
 wire \mem5_addr_b[2] ;
 wire \mem5_addr_b[3] ;
 wire \mem5_addr_b[4] ;
 wire \mem5_addr_b[5] ;
 wire \mem5_addr_b[6] ;
 wire \mem5_addr_b[7] ;
 wire \mem5_addr_b[8] ;
 wire \mem5_addr_b[9] ;
 wire mem5_cen_a;
 wire mem5_cen_b;
 wire mem5_clk_a;
 wire mem5_clk_b;
 wire \mem5_din_b[0] ;
 wire \mem5_din_b[10] ;
 wire \mem5_din_b[11] ;
 wire \mem5_din_b[12] ;
 wire \mem5_din_b[13] ;
 wire \mem5_din_b[14] ;
 wire \mem5_din_b[15] ;
 wire \mem5_din_b[16] ;
 wire \mem5_din_b[17] ;
 wire \mem5_din_b[18] ;
 wire \mem5_din_b[19] ;
 wire \mem5_din_b[1] ;
 wire \mem5_din_b[20] ;
 wire \mem5_din_b[21] ;
 wire \mem5_din_b[22] ;
 wire \mem5_din_b[23] ;
 wire \mem5_din_b[24] ;
 wire \mem5_din_b[25] ;
 wire \mem5_din_b[26] ;
 wire \mem5_din_b[27] ;
 wire \mem5_din_b[28] ;
 wire \mem5_din_b[29] ;
 wire \mem5_din_b[2] ;
 wire \mem5_din_b[30] ;
 wire \mem5_din_b[31] ;
 wire \mem5_din_b[3] ;
 wire \mem5_din_b[4] ;
 wire \mem5_din_b[5] ;
 wire \mem5_din_b[6] ;
 wire \mem5_din_b[7] ;
 wire \mem5_din_b[8] ;
 wire \mem5_din_b[9] ;
 wire \mem5_dout_a[0] ;
 wire \mem5_dout_a[10] ;
 wire \mem5_dout_a[11] ;
 wire \mem5_dout_a[12] ;
 wire \mem5_dout_a[13] ;
 wire \mem5_dout_a[14] ;
 wire \mem5_dout_a[15] ;
 wire \mem5_dout_a[16] ;
 wire \mem5_dout_a[17] ;
 wire \mem5_dout_a[18] ;
 wire \mem5_dout_a[19] ;
 wire \mem5_dout_a[1] ;
 wire \mem5_dout_a[20] ;
 wire \mem5_dout_a[21] ;
 wire \mem5_dout_a[22] ;
 wire \mem5_dout_a[23] ;
 wire \mem5_dout_a[24] ;
 wire \mem5_dout_a[25] ;
 wire \mem5_dout_a[26] ;
 wire \mem5_dout_a[27] ;
 wire \mem5_dout_a[28] ;
 wire \mem5_dout_a[29] ;
 wire \mem5_dout_a[2] ;
 wire \mem5_dout_a[30] ;
 wire \mem5_dout_a[31] ;
 wire \mem5_dout_a[3] ;
 wire \mem5_dout_a[4] ;
 wire \mem5_dout_a[5] ;
 wire \mem5_dout_a[6] ;
 wire \mem5_dout_a[7] ;
 wire \mem5_dout_a[8] ;
 wire \mem5_dout_a[9] ;
 wire \mem5_mask_b[0] ;
 wire \mem5_mask_b[1] ;
 wire \mem5_mask_b[2] ;
 wire \mem5_mask_b[3] ;
 wire mem5_web_b;
 wire \mem6_addr_a[2] ;
 wire \mem6_addr_a[3] ;
 wire \mem6_addr_a[4] ;
 wire \mem6_addr_a[5] ;
 wire \mem6_addr_a[6] ;
 wire \mem6_addr_a[7] ;
 wire \mem6_addr_a[8] ;
 wire \mem6_addr_a[9] ;
 wire \mem6_addr_b[2] ;
 wire \mem6_addr_b[3] ;
 wire \mem6_addr_b[4] ;
 wire \mem6_addr_b[5] ;
 wire \mem6_addr_b[6] ;
 wire \mem6_addr_b[7] ;
 wire \mem6_addr_b[8] ;
 wire \mem6_addr_b[9] ;
 wire mem6_cen_a;
 wire mem6_cen_b;
 wire mem6_clk_a;
 wire mem6_clk_b;
 wire \mem6_din_b[0] ;
 wire \mem6_din_b[10] ;
 wire \mem6_din_b[11] ;
 wire \mem6_din_b[12] ;
 wire \mem6_din_b[13] ;
 wire \mem6_din_b[14] ;
 wire \mem6_din_b[15] ;
 wire \mem6_din_b[16] ;
 wire \mem6_din_b[17] ;
 wire \mem6_din_b[18] ;
 wire \mem6_din_b[19] ;
 wire \mem6_din_b[1] ;
 wire \mem6_din_b[20] ;
 wire \mem6_din_b[21] ;
 wire \mem6_din_b[22] ;
 wire \mem6_din_b[23] ;
 wire \mem6_din_b[24] ;
 wire \mem6_din_b[25] ;
 wire \mem6_din_b[26] ;
 wire \mem6_din_b[27] ;
 wire \mem6_din_b[28] ;
 wire \mem6_din_b[29] ;
 wire \mem6_din_b[2] ;
 wire \mem6_din_b[30] ;
 wire \mem6_din_b[31] ;
 wire \mem6_din_b[3] ;
 wire \mem6_din_b[4] ;
 wire \mem6_din_b[5] ;
 wire \mem6_din_b[6] ;
 wire \mem6_din_b[7] ;
 wire \mem6_din_b[8] ;
 wire \mem6_din_b[9] ;
 wire \mem6_dout_a[0] ;
 wire \mem6_dout_a[10] ;
 wire \mem6_dout_a[11] ;
 wire \mem6_dout_a[12] ;
 wire \mem6_dout_a[13] ;
 wire \mem6_dout_a[14] ;
 wire \mem6_dout_a[15] ;
 wire \mem6_dout_a[16] ;
 wire \mem6_dout_a[17] ;
 wire \mem6_dout_a[18] ;
 wire \mem6_dout_a[19] ;
 wire \mem6_dout_a[1] ;
 wire \mem6_dout_a[20] ;
 wire \mem6_dout_a[21] ;
 wire \mem6_dout_a[22] ;
 wire \mem6_dout_a[23] ;
 wire \mem6_dout_a[24] ;
 wire \mem6_dout_a[25] ;
 wire \mem6_dout_a[26] ;
 wire \mem6_dout_a[27] ;
 wire \mem6_dout_a[28] ;
 wire \mem6_dout_a[29] ;
 wire \mem6_dout_a[2] ;
 wire \mem6_dout_a[30] ;
 wire \mem6_dout_a[31] ;
 wire \mem6_dout_a[3] ;
 wire \mem6_dout_a[4] ;
 wire \mem6_dout_a[5] ;
 wire \mem6_dout_a[6] ;
 wire \mem6_dout_a[7] ;
 wire \mem6_dout_a[8] ;
 wire \mem6_dout_a[9] ;
 wire \mem6_mask_b[0] ;
 wire \mem6_mask_b[1] ;
 wire \mem6_mask_b[2] ;
 wire \mem6_mask_b[3] ;
 wire mem6_web_b;
 wire \mem7_addr_a[2] ;
 wire \mem7_addr_a[3] ;
 wire \mem7_addr_a[4] ;
 wire \mem7_addr_a[5] ;
 wire \mem7_addr_a[6] ;
 wire \mem7_addr_a[7] ;
 wire \mem7_addr_a[8] ;
 wire \mem7_addr_a[9] ;
 wire \mem7_addr_b[2] ;
 wire \mem7_addr_b[3] ;
 wire \mem7_addr_b[4] ;
 wire \mem7_addr_b[5] ;
 wire \mem7_addr_b[6] ;
 wire \mem7_addr_b[7] ;
 wire \mem7_addr_b[8] ;
 wire \mem7_addr_b[9] ;
 wire mem7_cen_a;
 wire mem7_cen_b;
 wire mem7_clk_a;
 wire mem7_clk_b;
 wire \mem7_din_b[0] ;
 wire \mem7_din_b[10] ;
 wire \mem7_din_b[11] ;
 wire \mem7_din_b[12] ;
 wire \mem7_din_b[13] ;
 wire \mem7_din_b[14] ;
 wire \mem7_din_b[15] ;
 wire \mem7_din_b[16] ;
 wire \mem7_din_b[17] ;
 wire \mem7_din_b[18] ;
 wire \mem7_din_b[19] ;
 wire \mem7_din_b[1] ;
 wire \mem7_din_b[20] ;
 wire \mem7_din_b[21] ;
 wire \mem7_din_b[22] ;
 wire \mem7_din_b[23] ;
 wire \mem7_din_b[24] ;
 wire \mem7_din_b[25] ;
 wire \mem7_din_b[26] ;
 wire \mem7_din_b[27] ;
 wire \mem7_din_b[28] ;
 wire \mem7_din_b[29] ;
 wire \mem7_din_b[2] ;
 wire \mem7_din_b[30] ;
 wire \mem7_din_b[31] ;
 wire \mem7_din_b[3] ;
 wire \mem7_din_b[4] ;
 wire \mem7_din_b[5] ;
 wire \mem7_din_b[6] ;
 wire \mem7_din_b[7] ;
 wire \mem7_din_b[8] ;
 wire \mem7_din_b[9] ;
 wire \mem7_dout_a[0] ;
 wire \mem7_dout_a[10] ;
 wire \mem7_dout_a[11] ;
 wire \mem7_dout_a[12] ;
 wire \mem7_dout_a[13] ;
 wire \mem7_dout_a[14] ;
 wire \mem7_dout_a[15] ;
 wire \mem7_dout_a[16] ;
 wire \mem7_dout_a[17] ;
 wire \mem7_dout_a[18] ;
 wire \mem7_dout_a[19] ;
 wire \mem7_dout_a[1] ;
 wire \mem7_dout_a[20] ;
 wire \mem7_dout_a[21] ;
 wire \mem7_dout_a[22] ;
 wire \mem7_dout_a[23] ;
 wire \mem7_dout_a[24] ;
 wire \mem7_dout_a[25] ;
 wire \mem7_dout_a[26] ;
 wire \mem7_dout_a[27] ;
 wire \mem7_dout_a[28] ;
 wire \mem7_dout_a[29] ;
 wire \mem7_dout_a[2] ;
 wire \mem7_dout_a[30] ;
 wire \mem7_dout_a[31] ;
 wire \mem7_dout_a[3] ;
 wire \mem7_dout_a[4] ;
 wire \mem7_dout_a[5] ;
 wire \mem7_dout_a[6] ;
 wire \mem7_dout_a[7] ;
 wire \mem7_dout_a[8] ;
 wire \mem7_dout_a[9] ;
 wire \mem7_mask_b[0] ;
 wire \mem7_mask_b[1] ;
 wire \mem7_mask_b[2] ;
 wire \mem7_mask_b[3] ;
 wire mem7_web_b;
 wire \mem8_addr_a[2] ;
 wire \mem8_addr_a[3] ;
 wire \mem8_addr_a[4] ;
 wire \mem8_addr_a[5] ;
 wire \mem8_addr_a[6] ;
 wire \mem8_addr_a[7] ;
 wire \mem8_addr_a[8] ;
 wire \mem8_addr_a[9] ;
 wire \mem8_addr_b[2] ;
 wire \mem8_addr_b[3] ;
 wire \mem8_addr_b[4] ;
 wire \mem8_addr_b[5] ;
 wire \mem8_addr_b[6] ;
 wire \mem8_addr_b[7] ;
 wire \mem8_addr_b[8] ;
 wire \mem8_addr_b[9] ;
 wire mem8_cen_a;
 wire mem8_cen_b;
 wire mem8_clk_a;
 wire mem8_clk_b;
 wire \mem8_din_b[0] ;
 wire \mem8_din_b[10] ;
 wire \mem8_din_b[11] ;
 wire \mem8_din_b[12] ;
 wire \mem8_din_b[13] ;
 wire \mem8_din_b[14] ;
 wire \mem8_din_b[15] ;
 wire \mem8_din_b[16] ;
 wire \mem8_din_b[17] ;
 wire \mem8_din_b[18] ;
 wire \mem8_din_b[19] ;
 wire \mem8_din_b[1] ;
 wire \mem8_din_b[20] ;
 wire \mem8_din_b[21] ;
 wire \mem8_din_b[22] ;
 wire \mem8_din_b[23] ;
 wire \mem8_din_b[24] ;
 wire \mem8_din_b[25] ;
 wire \mem8_din_b[26] ;
 wire \mem8_din_b[27] ;
 wire \mem8_din_b[28] ;
 wire \mem8_din_b[29] ;
 wire \mem8_din_b[2] ;
 wire \mem8_din_b[30] ;
 wire \mem8_din_b[31] ;
 wire \mem8_din_b[3] ;
 wire \mem8_din_b[4] ;
 wire \mem8_din_b[5] ;
 wire \mem8_din_b[6] ;
 wire \mem8_din_b[7] ;
 wire \mem8_din_b[8] ;
 wire \mem8_din_b[9] ;
 wire \mem8_dout_a[0] ;
 wire \mem8_dout_a[10] ;
 wire \mem8_dout_a[11] ;
 wire \mem8_dout_a[12] ;
 wire \mem8_dout_a[13] ;
 wire \mem8_dout_a[14] ;
 wire \mem8_dout_a[15] ;
 wire \mem8_dout_a[16] ;
 wire \mem8_dout_a[17] ;
 wire \mem8_dout_a[18] ;
 wire \mem8_dout_a[19] ;
 wire \mem8_dout_a[1] ;
 wire \mem8_dout_a[20] ;
 wire \mem8_dout_a[21] ;
 wire \mem8_dout_a[22] ;
 wire \mem8_dout_a[23] ;
 wire \mem8_dout_a[24] ;
 wire \mem8_dout_a[25] ;
 wire \mem8_dout_a[26] ;
 wire \mem8_dout_a[27] ;
 wire \mem8_dout_a[28] ;
 wire \mem8_dout_a[29] ;
 wire \mem8_dout_a[2] ;
 wire \mem8_dout_a[30] ;
 wire \mem8_dout_a[31] ;
 wire \mem8_dout_a[3] ;
 wire \mem8_dout_a[4] ;
 wire \mem8_dout_a[5] ;
 wire \mem8_dout_a[6] ;
 wire \mem8_dout_a[7] ;
 wire \mem8_dout_a[8] ;
 wire \mem8_dout_a[9] ;
 wire \mem8_mask_b[0] ;
 wire \mem8_mask_b[1] ;
 wire \mem8_mask_b[2] ;
 wire \mem8_mask_b[3] ;
 wire mem8_web_b;
 wire scan_clk;
 wire scan_en;
 wire scan_en_glbl;
 wire scan_en_mbist1;
 wire scan_en_mbist2;
 wire scan_en_mbist3;
 wire scan_en_mbist4;
 wire scan_en_mbist5;
 wire scan_en_mbist6;
 wire scan_en_mbist7;
 wire scan_en_mbist8;
 wire scan_en_wbi;
 wire \scan_in[0] ;
 wire \scan_in[1] ;
 wire \scan_in[2] ;
 wire \scan_in[3] ;
 wire \scan_in[4] ;
 wire \scan_in[5] ;
 wire \scan_in[6] ;
 wire \scan_in[7] ;
 wire scan_mode;
 wire scan_mode_glbl;
 wire scan_mode_mbist1;
 wire scan_mode_mbist2;
 wire scan_mode_mbist3;
 wire scan_mode_mbist4;
 wire scan_mode_mbist5;
 wire scan_mode_mbist6;
 wire scan_mode_mbist7;
 wire scan_mode_mbist8;
 wire scan_mode_wbi;
 wire \scan_out_glbl[0] ;
 wire \scan_out_glbl[1] ;
 wire \scan_out_glbl[2] ;
 wire \scan_out_glbl[3] ;
 wire \scan_out_glbl[4] ;
 wire \scan_out_glbl[5] ;
 wire \scan_out_glbl[6] ;
 wire \scan_out_glbl[7] ;
 wire \scan_out_mbist1[0] ;
 wire \scan_out_mbist1[1] ;
 wire \scan_out_mbist1[2] ;
 wire \scan_out_mbist1[3] ;
 wire \scan_out_mbist1[4] ;
 wire \scan_out_mbist1[5] ;
 wire \scan_out_mbist1[6] ;
 wire \scan_out_mbist1[7] ;
 wire \scan_out_mbist2[0] ;
 wire \scan_out_mbist2[1] ;
 wire \scan_out_mbist2[2] ;
 wire \scan_out_mbist2[3] ;
 wire \scan_out_mbist2[4] ;
 wire \scan_out_mbist2[5] ;
 wire \scan_out_mbist2[6] ;
 wire \scan_out_mbist2[7] ;
 wire \scan_out_mbist3[0] ;
 wire \scan_out_mbist3[1] ;
 wire \scan_out_mbist3[2] ;
 wire \scan_out_mbist3[3] ;
 wire \scan_out_mbist3[4] ;
 wire \scan_out_mbist3[5] ;
 wire \scan_out_mbist3[6] ;
 wire \scan_out_mbist3[7] ;
 wire \scan_out_mbist4[0] ;
 wire \scan_out_mbist4[1] ;
 wire \scan_out_mbist4[2] ;
 wire \scan_out_mbist4[3] ;
 wire \scan_out_mbist4[4] ;
 wire \scan_out_mbist4[5] ;
 wire \scan_out_mbist4[6] ;
 wire \scan_out_mbist4[7] ;
 wire \scan_out_mbist5[0] ;
 wire \scan_out_mbist5[1] ;
 wire \scan_out_mbist5[2] ;
 wire \scan_out_mbist5[3] ;
 wire \scan_out_mbist5[4] ;
 wire \scan_out_mbist5[5] ;
 wire \scan_out_mbist5[6] ;
 wire \scan_out_mbist5[7] ;
 wire \scan_out_mbist6[0] ;
 wire \scan_out_mbist6[1] ;
 wire \scan_out_mbist6[2] ;
 wire \scan_out_mbist6[3] ;
 wire \scan_out_mbist6[4] ;
 wire \scan_out_mbist6[5] ;
 wire \scan_out_mbist6[6] ;
 wire \scan_out_mbist6[7] ;
 wire \scan_out_mbist7[0] ;
 wire \scan_out_mbist7[1] ;
 wire \scan_out_mbist7[2] ;
 wire \scan_out_mbist7[3] ;
 wire \scan_out_mbist7[4] ;
 wire \scan_out_mbist7[5] ;
 wire \scan_out_mbist7[6] ;
 wire \scan_out_mbist7[7] ;
 wire \scan_out_mbist8[0] ;
 wire \scan_out_mbist8[1] ;
 wire \scan_out_mbist8[2] ;
 wire \scan_out_mbist8[3] ;
 wire \scan_out_mbist8[4] ;
 wire \scan_out_mbist8[5] ;
 wire \scan_out_mbist8[6] ;
 wire \scan_out_mbist8[7] ;
 wire \scan_out_wbi[0] ;
 wire \scan_out_wbi[1] ;
 wire \scan_out_wbi[2] ;
 wire \scan_out_wbi[3] ;
 wire \scan_out_wbi[4] ;
 wire \scan_out_wbi[5] ;
 wire \scan_out_wbi[6] ;
 wire \scan_out_wbi[7] ;
 wire scan_rst_n;
 wire wbd_clk_glbl;
 wire wbd_clk_glbl_int;
 wire wbd_clk_int;
 wire wbd_clk_mbist1;
 wire wbd_clk_mbist1_int;
 wire wbd_clk_mbist2;
 wire wbd_clk_mbist2_int;
 wire wbd_clk_mbist3;
 wire wbd_clk_mbist3_int;
 wire wbd_clk_mbist4;
 wire wbd_clk_mbist4_int;
 wire wbd_clk_mbist5;
 wire wbd_clk_mbist5_int;
 wire wbd_clk_mbist6;
 wire wbd_clk_mbist6_int;
 wire wbd_clk_mbist7;
 wire wbd_clk_mbist7_int;
 wire wbd_clk_mbist8;
 wire wbd_clk_mbist8_int;
 wire wbd_clk_wh;
 wire wbd_clk_wi;
 wire wbd_glbl_ack_i;
 wire \wbd_glbl_adr_o[0] ;
 wire \wbd_glbl_adr_o[1] ;
 wire \wbd_glbl_adr_o[2] ;
 wire \wbd_glbl_adr_o[3] ;
 wire \wbd_glbl_adr_o[4] ;
 wire \wbd_glbl_adr_o[5] ;
 wire \wbd_glbl_adr_o[6] ;
 wire \wbd_glbl_adr_o[7] ;
 wire wbd_glbl_cyc_o;
 wire \wbd_glbl_dat_i[0] ;
 wire \wbd_glbl_dat_i[10] ;
 wire \wbd_glbl_dat_i[11] ;
 wire \wbd_glbl_dat_i[12] ;
 wire \wbd_glbl_dat_i[13] ;
 wire \wbd_glbl_dat_i[14] ;
 wire \wbd_glbl_dat_i[15] ;
 wire \wbd_glbl_dat_i[16] ;
 wire \wbd_glbl_dat_i[17] ;
 wire \wbd_glbl_dat_i[18] ;
 wire \wbd_glbl_dat_i[19] ;
 wire \wbd_glbl_dat_i[1] ;
 wire \wbd_glbl_dat_i[20] ;
 wire \wbd_glbl_dat_i[21] ;
 wire \wbd_glbl_dat_i[22] ;
 wire \wbd_glbl_dat_i[23] ;
 wire \wbd_glbl_dat_i[24] ;
 wire \wbd_glbl_dat_i[25] ;
 wire \wbd_glbl_dat_i[26] ;
 wire \wbd_glbl_dat_i[27] ;
 wire \wbd_glbl_dat_i[28] ;
 wire \wbd_glbl_dat_i[29] ;
 wire \wbd_glbl_dat_i[2] ;
 wire \wbd_glbl_dat_i[30] ;
 wire \wbd_glbl_dat_i[31] ;
 wire \wbd_glbl_dat_i[3] ;
 wire \wbd_glbl_dat_i[4] ;
 wire \wbd_glbl_dat_i[5] ;
 wire \wbd_glbl_dat_i[6] ;
 wire \wbd_glbl_dat_i[7] ;
 wire \wbd_glbl_dat_i[8] ;
 wire \wbd_glbl_dat_i[9] ;
 wire \wbd_glbl_dat_o[0] ;
 wire \wbd_glbl_dat_o[10] ;
 wire \wbd_glbl_dat_o[11] ;
 wire \wbd_glbl_dat_o[12] ;
 wire \wbd_glbl_dat_o[13] ;
 wire \wbd_glbl_dat_o[14] ;
 wire \wbd_glbl_dat_o[15] ;
 wire \wbd_glbl_dat_o[16] ;
 wire \wbd_glbl_dat_o[17] ;
 wire \wbd_glbl_dat_o[18] ;
 wire \wbd_glbl_dat_o[19] ;
 wire \wbd_glbl_dat_o[1] ;
 wire \wbd_glbl_dat_o[20] ;
 wire \wbd_glbl_dat_o[21] ;
 wire \wbd_glbl_dat_o[22] ;
 wire \wbd_glbl_dat_o[23] ;
 wire \wbd_glbl_dat_o[24] ;
 wire \wbd_glbl_dat_o[25] ;
 wire \wbd_glbl_dat_o[26] ;
 wire \wbd_glbl_dat_o[27] ;
 wire \wbd_glbl_dat_o[28] ;
 wire \wbd_glbl_dat_o[29] ;
 wire \wbd_glbl_dat_o[2] ;
 wire \wbd_glbl_dat_o[30] ;
 wire \wbd_glbl_dat_o[31] ;
 wire \wbd_glbl_dat_o[3] ;
 wire \wbd_glbl_dat_o[4] ;
 wire \wbd_glbl_dat_o[5] ;
 wire \wbd_glbl_dat_o[6] ;
 wire \wbd_glbl_dat_o[7] ;
 wire \wbd_glbl_dat_o[8] ;
 wire \wbd_glbl_dat_o[9] ;
 wire \wbd_glbl_sel_o[0] ;
 wire \wbd_glbl_sel_o[1] ;
 wire \wbd_glbl_sel_o[2] ;
 wire \wbd_glbl_sel_o[3] ;
 wire wbd_glbl_stb_o;
 wire wbd_glbl_we_o;
 wire wbd_int_ack_o;
 wire \wbd_int_adr_i[0] ;
 wire \wbd_int_adr_i[10] ;
 wire \wbd_int_adr_i[11] ;
 wire \wbd_int_adr_i[12] ;
 wire \wbd_int_adr_i[13] ;
 wire \wbd_int_adr_i[14] ;
 wire \wbd_int_adr_i[15] ;
 wire \wbd_int_adr_i[16] ;
 wire \wbd_int_adr_i[17] ;
 wire \wbd_int_adr_i[18] ;
 wire \wbd_int_adr_i[19] ;
 wire \wbd_int_adr_i[1] ;
 wire \wbd_int_adr_i[20] ;
 wire \wbd_int_adr_i[21] ;
 wire \wbd_int_adr_i[22] ;
 wire \wbd_int_adr_i[23] ;
 wire \wbd_int_adr_i[24] ;
 wire \wbd_int_adr_i[25] ;
 wire \wbd_int_adr_i[26] ;
 wire \wbd_int_adr_i[27] ;
 wire \wbd_int_adr_i[28] ;
 wire \wbd_int_adr_i[29] ;
 wire \wbd_int_adr_i[2] ;
 wire \wbd_int_adr_i[30] ;
 wire \wbd_int_adr_i[31] ;
 wire \wbd_int_adr_i[3] ;
 wire \wbd_int_adr_i[4] ;
 wire \wbd_int_adr_i[5] ;
 wire \wbd_int_adr_i[6] ;
 wire \wbd_int_adr_i[7] ;
 wire \wbd_int_adr_i[8] ;
 wire \wbd_int_adr_i[9] ;
 wire wbd_int_cyc_i;
 wire \wbd_int_dat_i[0] ;
 wire \wbd_int_dat_i[10] ;
 wire \wbd_int_dat_i[11] ;
 wire \wbd_int_dat_i[12] ;
 wire \wbd_int_dat_i[13] ;
 wire \wbd_int_dat_i[14] ;
 wire \wbd_int_dat_i[15] ;
 wire \wbd_int_dat_i[16] ;
 wire \wbd_int_dat_i[17] ;
 wire \wbd_int_dat_i[18] ;
 wire \wbd_int_dat_i[19] ;
 wire \wbd_int_dat_i[1] ;
 wire \wbd_int_dat_i[20] ;
 wire \wbd_int_dat_i[21] ;
 wire \wbd_int_dat_i[22] ;
 wire \wbd_int_dat_i[23] ;
 wire \wbd_int_dat_i[24] ;
 wire \wbd_int_dat_i[25] ;
 wire \wbd_int_dat_i[26] ;
 wire \wbd_int_dat_i[27] ;
 wire \wbd_int_dat_i[28] ;
 wire \wbd_int_dat_i[29] ;
 wire \wbd_int_dat_i[2] ;
 wire \wbd_int_dat_i[30] ;
 wire \wbd_int_dat_i[31] ;
 wire \wbd_int_dat_i[3] ;
 wire \wbd_int_dat_i[4] ;
 wire \wbd_int_dat_i[5] ;
 wire \wbd_int_dat_i[6] ;
 wire \wbd_int_dat_i[7] ;
 wire \wbd_int_dat_i[8] ;
 wire \wbd_int_dat_i[9] ;
 wire \wbd_int_dat_o[0] ;
 wire \wbd_int_dat_o[10] ;
 wire \wbd_int_dat_o[11] ;
 wire \wbd_int_dat_o[12] ;
 wire \wbd_int_dat_o[13] ;
 wire \wbd_int_dat_o[14] ;
 wire \wbd_int_dat_o[15] ;
 wire \wbd_int_dat_o[16] ;
 wire \wbd_int_dat_o[17] ;
 wire \wbd_int_dat_o[18] ;
 wire \wbd_int_dat_o[19] ;
 wire \wbd_int_dat_o[1] ;
 wire \wbd_int_dat_o[20] ;
 wire \wbd_int_dat_o[21] ;
 wire \wbd_int_dat_o[22] ;
 wire \wbd_int_dat_o[23] ;
 wire \wbd_int_dat_o[24] ;
 wire \wbd_int_dat_o[25] ;
 wire \wbd_int_dat_o[26] ;
 wire \wbd_int_dat_o[27] ;
 wire \wbd_int_dat_o[28] ;
 wire \wbd_int_dat_o[29] ;
 wire \wbd_int_dat_o[2] ;
 wire \wbd_int_dat_o[30] ;
 wire \wbd_int_dat_o[31] ;
 wire \wbd_int_dat_o[3] ;
 wire \wbd_int_dat_o[4] ;
 wire \wbd_int_dat_o[5] ;
 wire \wbd_int_dat_o[6] ;
 wire \wbd_int_dat_o[7] ;
 wire \wbd_int_dat_o[8] ;
 wire \wbd_int_dat_o[9] ;
 wire wbd_int_err_o;
 wire wbd_int_rst_n;
 wire \wbd_int_sel_i[0] ;
 wire \wbd_int_sel_i[1] ;
 wire \wbd_int_sel_i[2] ;
 wire \wbd_int_sel_i[3] ;
 wire wbd_int_stb_i;
 wire wbd_int_we_i;
 wire wbd_mbist1_ack_i;
 wire \wbd_mbist1_adr_o[0] ;
 wire \wbd_mbist1_adr_o[10] ;
 wire \wbd_mbist1_adr_o[1] ;
 wire \wbd_mbist1_adr_o[2] ;
 wire \wbd_mbist1_adr_o[3] ;
 wire \wbd_mbist1_adr_o[4] ;
 wire \wbd_mbist1_adr_o[5] ;
 wire \wbd_mbist1_adr_o[6] ;
 wire \wbd_mbist1_adr_o[7] ;
 wire \wbd_mbist1_adr_o[8] ;
 wire \wbd_mbist1_adr_o[9] ;
 wire wbd_mbist1_cyc_o;
 wire \wbd_mbist1_dat_i[0] ;
 wire \wbd_mbist1_dat_i[10] ;
 wire \wbd_mbist1_dat_i[11] ;
 wire \wbd_mbist1_dat_i[12] ;
 wire \wbd_mbist1_dat_i[13] ;
 wire \wbd_mbist1_dat_i[14] ;
 wire \wbd_mbist1_dat_i[15] ;
 wire \wbd_mbist1_dat_i[16] ;
 wire \wbd_mbist1_dat_i[17] ;
 wire \wbd_mbist1_dat_i[18] ;
 wire \wbd_mbist1_dat_i[19] ;
 wire \wbd_mbist1_dat_i[1] ;
 wire \wbd_mbist1_dat_i[20] ;
 wire \wbd_mbist1_dat_i[21] ;
 wire \wbd_mbist1_dat_i[22] ;
 wire \wbd_mbist1_dat_i[23] ;
 wire \wbd_mbist1_dat_i[24] ;
 wire \wbd_mbist1_dat_i[25] ;
 wire \wbd_mbist1_dat_i[26] ;
 wire \wbd_mbist1_dat_i[27] ;
 wire \wbd_mbist1_dat_i[28] ;
 wire \wbd_mbist1_dat_i[29] ;
 wire \wbd_mbist1_dat_i[2] ;
 wire \wbd_mbist1_dat_i[30] ;
 wire \wbd_mbist1_dat_i[31] ;
 wire \wbd_mbist1_dat_i[3] ;
 wire \wbd_mbist1_dat_i[4] ;
 wire \wbd_mbist1_dat_i[5] ;
 wire \wbd_mbist1_dat_i[6] ;
 wire \wbd_mbist1_dat_i[7] ;
 wire \wbd_mbist1_dat_i[8] ;
 wire \wbd_mbist1_dat_i[9] ;
 wire \wbd_mbist1_dat_o[0] ;
 wire \wbd_mbist1_dat_o[10] ;
 wire \wbd_mbist1_dat_o[11] ;
 wire \wbd_mbist1_dat_o[12] ;
 wire \wbd_mbist1_dat_o[13] ;
 wire \wbd_mbist1_dat_o[14] ;
 wire \wbd_mbist1_dat_o[15] ;
 wire \wbd_mbist1_dat_o[16] ;
 wire \wbd_mbist1_dat_o[17] ;
 wire \wbd_mbist1_dat_o[18] ;
 wire \wbd_mbist1_dat_o[19] ;
 wire \wbd_mbist1_dat_o[1] ;
 wire \wbd_mbist1_dat_o[20] ;
 wire \wbd_mbist1_dat_o[21] ;
 wire \wbd_mbist1_dat_o[22] ;
 wire \wbd_mbist1_dat_o[23] ;
 wire \wbd_mbist1_dat_o[24] ;
 wire \wbd_mbist1_dat_o[25] ;
 wire \wbd_mbist1_dat_o[26] ;
 wire \wbd_mbist1_dat_o[27] ;
 wire \wbd_mbist1_dat_o[28] ;
 wire \wbd_mbist1_dat_o[29] ;
 wire \wbd_mbist1_dat_o[2] ;
 wire \wbd_mbist1_dat_o[30] ;
 wire \wbd_mbist1_dat_o[31] ;
 wire \wbd_mbist1_dat_o[3] ;
 wire \wbd_mbist1_dat_o[4] ;
 wire \wbd_mbist1_dat_o[5] ;
 wire \wbd_mbist1_dat_o[6] ;
 wire \wbd_mbist1_dat_o[7] ;
 wire \wbd_mbist1_dat_o[8] ;
 wire \wbd_mbist1_dat_o[9] ;
 wire \wbd_mbist1_sel_o[0] ;
 wire \wbd_mbist1_sel_o[1] ;
 wire \wbd_mbist1_sel_o[2] ;
 wire \wbd_mbist1_sel_o[3] ;
 wire wbd_mbist1_stb_o;
 wire wbd_mbist1_we_o;
 wire wbd_mbist2_ack_i;
 wire \wbd_mbist2_adr_o[0] ;
 wire \wbd_mbist2_adr_o[10] ;
 wire \wbd_mbist2_adr_o[1] ;
 wire \wbd_mbist2_adr_o[2] ;
 wire \wbd_mbist2_adr_o[3] ;
 wire \wbd_mbist2_adr_o[4] ;
 wire \wbd_mbist2_adr_o[5] ;
 wire \wbd_mbist2_adr_o[6] ;
 wire \wbd_mbist2_adr_o[7] ;
 wire \wbd_mbist2_adr_o[8] ;
 wire \wbd_mbist2_adr_o[9] ;
 wire wbd_mbist2_cyc_o;
 wire \wbd_mbist2_dat_i[0] ;
 wire \wbd_mbist2_dat_i[10] ;
 wire \wbd_mbist2_dat_i[11] ;
 wire \wbd_mbist2_dat_i[12] ;
 wire \wbd_mbist2_dat_i[13] ;
 wire \wbd_mbist2_dat_i[14] ;
 wire \wbd_mbist2_dat_i[15] ;
 wire \wbd_mbist2_dat_i[16] ;
 wire \wbd_mbist2_dat_i[17] ;
 wire \wbd_mbist2_dat_i[18] ;
 wire \wbd_mbist2_dat_i[19] ;
 wire \wbd_mbist2_dat_i[1] ;
 wire \wbd_mbist2_dat_i[20] ;
 wire \wbd_mbist2_dat_i[21] ;
 wire \wbd_mbist2_dat_i[22] ;
 wire \wbd_mbist2_dat_i[23] ;
 wire \wbd_mbist2_dat_i[24] ;
 wire \wbd_mbist2_dat_i[25] ;
 wire \wbd_mbist2_dat_i[26] ;
 wire \wbd_mbist2_dat_i[27] ;
 wire \wbd_mbist2_dat_i[28] ;
 wire \wbd_mbist2_dat_i[29] ;
 wire \wbd_mbist2_dat_i[2] ;
 wire \wbd_mbist2_dat_i[30] ;
 wire \wbd_mbist2_dat_i[31] ;
 wire \wbd_mbist2_dat_i[3] ;
 wire \wbd_mbist2_dat_i[4] ;
 wire \wbd_mbist2_dat_i[5] ;
 wire \wbd_mbist2_dat_i[6] ;
 wire \wbd_mbist2_dat_i[7] ;
 wire \wbd_mbist2_dat_i[8] ;
 wire \wbd_mbist2_dat_i[9] ;
 wire \wbd_mbist2_dat_o[0] ;
 wire \wbd_mbist2_dat_o[10] ;
 wire \wbd_mbist2_dat_o[11] ;
 wire \wbd_mbist2_dat_o[12] ;
 wire \wbd_mbist2_dat_o[13] ;
 wire \wbd_mbist2_dat_o[14] ;
 wire \wbd_mbist2_dat_o[15] ;
 wire \wbd_mbist2_dat_o[16] ;
 wire \wbd_mbist2_dat_o[17] ;
 wire \wbd_mbist2_dat_o[18] ;
 wire \wbd_mbist2_dat_o[19] ;
 wire \wbd_mbist2_dat_o[1] ;
 wire \wbd_mbist2_dat_o[20] ;
 wire \wbd_mbist2_dat_o[21] ;
 wire \wbd_mbist2_dat_o[22] ;
 wire \wbd_mbist2_dat_o[23] ;
 wire \wbd_mbist2_dat_o[24] ;
 wire \wbd_mbist2_dat_o[25] ;
 wire \wbd_mbist2_dat_o[26] ;
 wire \wbd_mbist2_dat_o[27] ;
 wire \wbd_mbist2_dat_o[28] ;
 wire \wbd_mbist2_dat_o[29] ;
 wire \wbd_mbist2_dat_o[2] ;
 wire \wbd_mbist2_dat_o[30] ;
 wire \wbd_mbist2_dat_o[31] ;
 wire \wbd_mbist2_dat_o[3] ;
 wire \wbd_mbist2_dat_o[4] ;
 wire \wbd_mbist2_dat_o[5] ;
 wire \wbd_mbist2_dat_o[6] ;
 wire \wbd_mbist2_dat_o[7] ;
 wire \wbd_mbist2_dat_o[8] ;
 wire \wbd_mbist2_dat_o[9] ;
 wire \wbd_mbist2_sel_o[0] ;
 wire \wbd_mbist2_sel_o[1] ;
 wire \wbd_mbist2_sel_o[2] ;
 wire \wbd_mbist2_sel_o[3] ;
 wire wbd_mbist2_stb_o;
 wire wbd_mbist2_we_o;
 wire wbd_mbist3_ack_i;
 wire \wbd_mbist3_adr_o[0] ;
 wire \wbd_mbist3_adr_o[10] ;
 wire \wbd_mbist3_adr_o[1] ;
 wire \wbd_mbist3_adr_o[2] ;
 wire \wbd_mbist3_adr_o[3] ;
 wire \wbd_mbist3_adr_o[4] ;
 wire \wbd_mbist3_adr_o[5] ;
 wire \wbd_mbist3_adr_o[6] ;
 wire \wbd_mbist3_adr_o[7] ;
 wire \wbd_mbist3_adr_o[8] ;
 wire \wbd_mbist3_adr_o[9] ;
 wire wbd_mbist3_cyc_o;
 wire \wbd_mbist3_dat_i[0] ;
 wire \wbd_mbist3_dat_i[10] ;
 wire \wbd_mbist3_dat_i[11] ;
 wire \wbd_mbist3_dat_i[12] ;
 wire \wbd_mbist3_dat_i[13] ;
 wire \wbd_mbist3_dat_i[14] ;
 wire \wbd_mbist3_dat_i[15] ;
 wire \wbd_mbist3_dat_i[16] ;
 wire \wbd_mbist3_dat_i[17] ;
 wire \wbd_mbist3_dat_i[18] ;
 wire \wbd_mbist3_dat_i[19] ;
 wire \wbd_mbist3_dat_i[1] ;
 wire \wbd_mbist3_dat_i[20] ;
 wire \wbd_mbist3_dat_i[21] ;
 wire \wbd_mbist3_dat_i[22] ;
 wire \wbd_mbist3_dat_i[23] ;
 wire \wbd_mbist3_dat_i[24] ;
 wire \wbd_mbist3_dat_i[25] ;
 wire \wbd_mbist3_dat_i[26] ;
 wire \wbd_mbist3_dat_i[27] ;
 wire \wbd_mbist3_dat_i[28] ;
 wire \wbd_mbist3_dat_i[29] ;
 wire \wbd_mbist3_dat_i[2] ;
 wire \wbd_mbist3_dat_i[30] ;
 wire \wbd_mbist3_dat_i[31] ;
 wire \wbd_mbist3_dat_i[3] ;
 wire \wbd_mbist3_dat_i[4] ;
 wire \wbd_mbist3_dat_i[5] ;
 wire \wbd_mbist3_dat_i[6] ;
 wire \wbd_mbist3_dat_i[7] ;
 wire \wbd_mbist3_dat_i[8] ;
 wire \wbd_mbist3_dat_i[9] ;
 wire \wbd_mbist3_dat_o[0] ;
 wire \wbd_mbist3_dat_o[10] ;
 wire \wbd_mbist3_dat_o[11] ;
 wire \wbd_mbist3_dat_o[12] ;
 wire \wbd_mbist3_dat_o[13] ;
 wire \wbd_mbist3_dat_o[14] ;
 wire \wbd_mbist3_dat_o[15] ;
 wire \wbd_mbist3_dat_o[16] ;
 wire \wbd_mbist3_dat_o[17] ;
 wire \wbd_mbist3_dat_o[18] ;
 wire \wbd_mbist3_dat_o[19] ;
 wire \wbd_mbist3_dat_o[1] ;
 wire \wbd_mbist3_dat_o[20] ;
 wire \wbd_mbist3_dat_o[21] ;
 wire \wbd_mbist3_dat_o[22] ;
 wire \wbd_mbist3_dat_o[23] ;
 wire \wbd_mbist3_dat_o[24] ;
 wire \wbd_mbist3_dat_o[25] ;
 wire \wbd_mbist3_dat_o[26] ;
 wire \wbd_mbist3_dat_o[27] ;
 wire \wbd_mbist3_dat_o[28] ;
 wire \wbd_mbist3_dat_o[29] ;
 wire \wbd_mbist3_dat_o[2] ;
 wire \wbd_mbist3_dat_o[30] ;
 wire \wbd_mbist3_dat_o[31] ;
 wire \wbd_mbist3_dat_o[3] ;
 wire \wbd_mbist3_dat_o[4] ;
 wire \wbd_mbist3_dat_o[5] ;
 wire \wbd_mbist3_dat_o[6] ;
 wire \wbd_mbist3_dat_o[7] ;
 wire \wbd_mbist3_dat_o[8] ;
 wire \wbd_mbist3_dat_o[9] ;
 wire \wbd_mbist3_sel_o[0] ;
 wire \wbd_mbist3_sel_o[1] ;
 wire \wbd_mbist3_sel_o[2] ;
 wire \wbd_mbist3_sel_o[3] ;
 wire wbd_mbist3_stb_o;
 wire wbd_mbist3_we_o;
 wire wbd_mbist4_ack_i;
 wire \wbd_mbist4_adr_o[0] ;
 wire \wbd_mbist4_adr_o[10] ;
 wire \wbd_mbist4_adr_o[1] ;
 wire \wbd_mbist4_adr_o[2] ;
 wire \wbd_mbist4_adr_o[3] ;
 wire \wbd_mbist4_adr_o[4] ;
 wire \wbd_mbist4_adr_o[5] ;
 wire \wbd_mbist4_adr_o[6] ;
 wire \wbd_mbist4_adr_o[7] ;
 wire \wbd_mbist4_adr_o[8] ;
 wire \wbd_mbist4_adr_o[9] ;
 wire wbd_mbist4_cyc_o;
 wire \wbd_mbist4_dat_i[0] ;
 wire \wbd_mbist4_dat_i[10] ;
 wire \wbd_mbist4_dat_i[11] ;
 wire \wbd_mbist4_dat_i[12] ;
 wire \wbd_mbist4_dat_i[13] ;
 wire \wbd_mbist4_dat_i[14] ;
 wire \wbd_mbist4_dat_i[15] ;
 wire \wbd_mbist4_dat_i[16] ;
 wire \wbd_mbist4_dat_i[17] ;
 wire \wbd_mbist4_dat_i[18] ;
 wire \wbd_mbist4_dat_i[19] ;
 wire \wbd_mbist4_dat_i[1] ;
 wire \wbd_mbist4_dat_i[20] ;
 wire \wbd_mbist4_dat_i[21] ;
 wire \wbd_mbist4_dat_i[22] ;
 wire \wbd_mbist4_dat_i[23] ;
 wire \wbd_mbist4_dat_i[24] ;
 wire \wbd_mbist4_dat_i[25] ;
 wire \wbd_mbist4_dat_i[26] ;
 wire \wbd_mbist4_dat_i[27] ;
 wire \wbd_mbist4_dat_i[28] ;
 wire \wbd_mbist4_dat_i[29] ;
 wire \wbd_mbist4_dat_i[2] ;
 wire \wbd_mbist4_dat_i[30] ;
 wire \wbd_mbist4_dat_i[31] ;
 wire \wbd_mbist4_dat_i[3] ;
 wire \wbd_mbist4_dat_i[4] ;
 wire \wbd_mbist4_dat_i[5] ;
 wire \wbd_mbist4_dat_i[6] ;
 wire \wbd_mbist4_dat_i[7] ;
 wire \wbd_mbist4_dat_i[8] ;
 wire \wbd_mbist4_dat_i[9] ;
 wire \wbd_mbist4_dat_o[0] ;
 wire \wbd_mbist4_dat_o[10] ;
 wire \wbd_mbist4_dat_o[11] ;
 wire \wbd_mbist4_dat_o[12] ;
 wire \wbd_mbist4_dat_o[13] ;
 wire \wbd_mbist4_dat_o[14] ;
 wire \wbd_mbist4_dat_o[15] ;
 wire \wbd_mbist4_dat_o[16] ;
 wire \wbd_mbist4_dat_o[17] ;
 wire \wbd_mbist4_dat_o[18] ;
 wire \wbd_mbist4_dat_o[19] ;
 wire \wbd_mbist4_dat_o[1] ;
 wire \wbd_mbist4_dat_o[20] ;
 wire \wbd_mbist4_dat_o[21] ;
 wire \wbd_mbist4_dat_o[22] ;
 wire \wbd_mbist4_dat_o[23] ;
 wire \wbd_mbist4_dat_o[24] ;
 wire \wbd_mbist4_dat_o[25] ;
 wire \wbd_mbist4_dat_o[26] ;
 wire \wbd_mbist4_dat_o[27] ;
 wire \wbd_mbist4_dat_o[28] ;
 wire \wbd_mbist4_dat_o[29] ;
 wire \wbd_mbist4_dat_o[2] ;
 wire \wbd_mbist4_dat_o[30] ;
 wire \wbd_mbist4_dat_o[31] ;
 wire \wbd_mbist4_dat_o[3] ;
 wire \wbd_mbist4_dat_o[4] ;
 wire \wbd_mbist4_dat_o[5] ;
 wire \wbd_mbist4_dat_o[6] ;
 wire \wbd_mbist4_dat_o[7] ;
 wire \wbd_mbist4_dat_o[8] ;
 wire \wbd_mbist4_dat_o[9] ;
 wire \wbd_mbist4_sel_o[0] ;
 wire \wbd_mbist4_sel_o[1] ;
 wire \wbd_mbist4_sel_o[2] ;
 wire \wbd_mbist4_sel_o[3] ;
 wire wbd_mbist4_stb_o;
 wire wbd_mbist4_we_o;
 wire wbd_mbist5_ack_i;
 wire \wbd_mbist5_adr_o[0] ;
 wire \wbd_mbist5_adr_o[1] ;
 wire \wbd_mbist5_adr_o[2] ;
 wire \wbd_mbist5_adr_o[3] ;
 wire \wbd_mbist5_adr_o[4] ;
 wire \wbd_mbist5_adr_o[5] ;
 wire \wbd_mbist5_adr_o[6] ;
 wire \wbd_mbist5_adr_o[7] ;
 wire \wbd_mbist5_adr_o[8] ;
 wire \wbd_mbist5_adr_o[9] ;
 wire wbd_mbist5_cyc_o;
 wire \wbd_mbist5_dat_i[0] ;
 wire \wbd_mbist5_dat_i[10] ;
 wire \wbd_mbist5_dat_i[11] ;
 wire \wbd_mbist5_dat_i[12] ;
 wire \wbd_mbist5_dat_i[13] ;
 wire \wbd_mbist5_dat_i[14] ;
 wire \wbd_mbist5_dat_i[15] ;
 wire \wbd_mbist5_dat_i[16] ;
 wire \wbd_mbist5_dat_i[17] ;
 wire \wbd_mbist5_dat_i[18] ;
 wire \wbd_mbist5_dat_i[19] ;
 wire \wbd_mbist5_dat_i[1] ;
 wire \wbd_mbist5_dat_i[20] ;
 wire \wbd_mbist5_dat_i[21] ;
 wire \wbd_mbist5_dat_i[22] ;
 wire \wbd_mbist5_dat_i[23] ;
 wire \wbd_mbist5_dat_i[24] ;
 wire \wbd_mbist5_dat_i[25] ;
 wire \wbd_mbist5_dat_i[26] ;
 wire \wbd_mbist5_dat_i[27] ;
 wire \wbd_mbist5_dat_i[28] ;
 wire \wbd_mbist5_dat_i[29] ;
 wire \wbd_mbist5_dat_i[2] ;
 wire \wbd_mbist5_dat_i[30] ;
 wire \wbd_mbist5_dat_i[31] ;
 wire \wbd_mbist5_dat_i[3] ;
 wire \wbd_mbist5_dat_i[4] ;
 wire \wbd_mbist5_dat_i[5] ;
 wire \wbd_mbist5_dat_i[6] ;
 wire \wbd_mbist5_dat_i[7] ;
 wire \wbd_mbist5_dat_i[8] ;
 wire \wbd_mbist5_dat_i[9] ;
 wire \wbd_mbist5_dat_o[0] ;
 wire \wbd_mbist5_dat_o[10] ;
 wire \wbd_mbist5_dat_o[11] ;
 wire \wbd_mbist5_dat_o[12] ;
 wire \wbd_mbist5_dat_o[13] ;
 wire \wbd_mbist5_dat_o[14] ;
 wire \wbd_mbist5_dat_o[15] ;
 wire \wbd_mbist5_dat_o[16] ;
 wire \wbd_mbist5_dat_o[17] ;
 wire \wbd_mbist5_dat_o[18] ;
 wire \wbd_mbist5_dat_o[19] ;
 wire \wbd_mbist5_dat_o[1] ;
 wire \wbd_mbist5_dat_o[20] ;
 wire \wbd_mbist5_dat_o[21] ;
 wire \wbd_mbist5_dat_o[22] ;
 wire \wbd_mbist5_dat_o[23] ;
 wire \wbd_mbist5_dat_o[24] ;
 wire \wbd_mbist5_dat_o[25] ;
 wire \wbd_mbist5_dat_o[26] ;
 wire \wbd_mbist5_dat_o[27] ;
 wire \wbd_mbist5_dat_o[28] ;
 wire \wbd_mbist5_dat_o[29] ;
 wire \wbd_mbist5_dat_o[2] ;
 wire \wbd_mbist5_dat_o[30] ;
 wire \wbd_mbist5_dat_o[31] ;
 wire \wbd_mbist5_dat_o[3] ;
 wire \wbd_mbist5_dat_o[4] ;
 wire \wbd_mbist5_dat_o[5] ;
 wire \wbd_mbist5_dat_o[6] ;
 wire \wbd_mbist5_dat_o[7] ;
 wire \wbd_mbist5_dat_o[8] ;
 wire \wbd_mbist5_dat_o[9] ;
 wire \wbd_mbist5_sel_o[0] ;
 wire \wbd_mbist5_sel_o[1] ;
 wire \wbd_mbist5_sel_o[2] ;
 wire \wbd_mbist5_sel_o[3] ;
 wire wbd_mbist5_stb_o;
 wire wbd_mbist5_we_o;
 wire wbd_mbist6_ack_i;
 wire \wbd_mbist6_adr_o[0] ;
 wire \wbd_mbist6_adr_o[1] ;
 wire \wbd_mbist6_adr_o[2] ;
 wire \wbd_mbist6_adr_o[3] ;
 wire \wbd_mbist6_adr_o[4] ;
 wire \wbd_mbist6_adr_o[5] ;
 wire \wbd_mbist6_adr_o[6] ;
 wire \wbd_mbist6_adr_o[7] ;
 wire \wbd_mbist6_adr_o[8] ;
 wire \wbd_mbist6_adr_o[9] ;
 wire wbd_mbist6_cyc_o;
 wire \wbd_mbist6_dat_i[0] ;
 wire \wbd_mbist6_dat_i[10] ;
 wire \wbd_mbist6_dat_i[11] ;
 wire \wbd_mbist6_dat_i[12] ;
 wire \wbd_mbist6_dat_i[13] ;
 wire \wbd_mbist6_dat_i[14] ;
 wire \wbd_mbist6_dat_i[15] ;
 wire \wbd_mbist6_dat_i[16] ;
 wire \wbd_mbist6_dat_i[17] ;
 wire \wbd_mbist6_dat_i[18] ;
 wire \wbd_mbist6_dat_i[19] ;
 wire \wbd_mbist6_dat_i[1] ;
 wire \wbd_mbist6_dat_i[20] ;
 wire \wbd_mbist6_dat_i[21] ;
 wire \wbd_mbist6_dat_i[22] ;
 wire \wbd_mbist6_dat_i[23] ;
 wire \wbd_mbist6_dat_i[24] ;
 wire \wbd_mbist6_dat_i[25] ;
 wire \wbd_mbist6_dat_i[26] ;
 wire \wbd_mbist6_dat_i[27] ;
 wire \wbd_mbist6_dat_i[28] ;
 wire \wbd_mbist6_dat_i[29] ;
 wire \wbd_mbist6_dat_i[2] ;
 wire \wbd_mbist6_dat_i[30] ;
 wire \wbd_mbist6_dat_i[31] ;
 wire \wbd_mbist6_dat_i[3] ;
 wire \wbd_mbist6_dat_i[4] ;
 wire \wbd_mbist6_dat_i[5] ;
 wire \wbd_mbist6_dat_i[6] ;
 wire \wbd_mbist6_dat_i[7] ;
 wire \wbd_mbist6_dat_i[8] ;
 wire \wbd_mbist6_dat_i[9] ;
 wire \wbd_mbist6_dat_o[0] ;
 wire \wbd_mbist6_dat_o[10] ;
 wire \wbd_mbist6_dat_o[11] ;
 wire \wbd_mbist6_dat_o[12] ;
 wire \wbd_mbist6_dat_o[13] ;
 wire \wbd_mbist6_dat_o[14] ;
 wire \wbd_mbist6_dat_o[15] ;
 wire \wbd_mbist6_dat_o[16] ;
 wire \wbd_mbist6_dat_o[17] ;
 wire \wbd_mbist6_dat_o[18] ;
 wire \wbd_mbist6_dat_o[19] ;
 wire \wbd_mbist6_dat_o[1] ;
 wire \wbd_mbist6_dat_o[20] ;
 wire \wbd_mbist6_dat_o[21] ;
 wire \wbd_mbist6_dat_o[22] ;
 wire \wbd_mbist6_dat_o[23] ;
 wire \wbd_mbist6_dat_o[24] ;
 wire \wbd_mbist6_dat_o[25] ;
 wire \wbd_mbist6_dat_o[26] ;
 wire \wbd_mbist6_dat_o[27] ;
 wire \wbd_mbist6_dat_o[28] ;
 wire \wbd_mbist6_dat_o[29] ;
 wire \wbd_mbist6_dat_o[2] ;
 wire \wbd_mbist6_dat_o[30] ;
 wire \wbd_mbist6_dat_o[31] ;
 wire \wbd_mbist6_dat_o[3] ;
 wire \wbd_mbist6_dat_o[4] ;
 wire \wbd_mbist6_dat_o[5] ;
 wire \wbd_mbist6_dat_o[6] ;
 wire \wbd_mbist6_dat_o[7] ;
 wire \wbd_mbist6_dat_o[8] ;
 wire \wbd_mbist6_dat_o[9] ;
 wire \wbd_mbist6_sel_o[0] ;
 wire \wbd_mbist6_sel_o[1] ;
 wire \wbd_mbist6_sel_o[2] ;
 wire \wbd_mbist6_sel_o[3] ;
 wire wbd_mbist6_stb_o;
 wire wbd_mbist6_we_o;
 wire wbd_mbist7_ack_i;
 wire \wbd_mbist7_adr_o[0] ;
 wire \wbd_mbist7_adr_o[1] ;
 wire \wbd_mbist7_adr_o[2] ;
 wire \wbd_mbist7_adr_o[3] ;
 wire \wbd_mbist7_adr_o[4] ;
 wire \wbd_mbist7_adr_o[5] ;
 wire \wbd_mbist7_adr_o[6] ;
 wire \wbd_mbist7_adr_o[7] ;
 wire \wbd_mbist7_adr_o[8] ;
 wire \wbd_mbist7_adr_o[9] ;
 wire wbd_mbist7_cyc_o;
 wire \wbd_mbist7_dat_i[0] ;
 wire \wbd_mbist7_dat_i[10] ;
 wire \wbd_mbist7_dat_i[11] ;
 wire \wbd_mbist7_dat_i[12] ;
 wire \wbd_mbist7_dat_i[13] ;
 wire \wbd_mbist7_dat_i[14] ;
 wire \wbd_mbist7_dat_i[15] ;
 wire \wbd_mbist7_dat_i[16] ;
 wire \wbd_mbist7_dat_i[17] ;
 wire \wbd_mbist7_dat_i[18] ;
 wire \wbd_mbist7_dat_i[19] ;
 wire \wbd_mbist7_dat_i[1] ;
 wire \wbd_mbist7_dat_i[20] ;
 wire \wbd_mbist7_dat_i[21] ;
 wire \wbd_mbist7_dat_i[22] ;
 wire \wbd_mbist7_dat_i[23] ;
 wire \wbd_mbist7_dat_i[24] ;
 wire \wbd_mbist7_dat_i[25] ;
 wire \wbd_mbist7_dat_i[26] ;
 wire \wbd_mbist7_dat_i[27] ;
 wire \wbd_mbist7_dat_i[28] ;
 wire \wbd_mbist7_dat_i[29] ;
 wire \wbd_mbist7_dat_i[2] ;
 wire \wbd_mbist7_dat_i[30] ;
 wire \wbd_mbist7_dat_i[31] ;
 wire \wbd_mbist7_dat_i[3] ;
 wire \wbd_mbist7_dat_i[4] ;
 wire \wbd_mbist7_dat_i[5] ;
 wire \wbd_mbist7_dat_i[6] ;
 wire \wbd_mbist7_dat_i[7] ;
 wire \wbd_mbist7_dat_i[8] ;
 wire \wbd_mbist7_dat_i[9] ;
 wire \wbd_mbist7_dat_o[0] ;
 wire \wbd_mbist7_dat_o[10] ;
 wire \wbd_mbist7_dat_o[11] ;
 wire \wbd_mbist7_dat_o[12] ;
 wire \wbd_mbist7_dat_o[13] ;
 wire \wbd_mbist7_dat_o[14] ;
 wire \wbd_mbist7_dat_o[15] ;
 wire \wbd_mbist7_dat_o[16] ;
 wire \wbd_mbist7_dat_o[17] ;
 wire \wbd_mbist7_dat_o[18] ;
 wire \wbd_mbist7_dat_o[19] ;
 wire \wbd_mbist7_dat_o[1] ;
 wire \wbd_mbist7_dat_o[20] ;
 wire \wbd_mbist7_dat_o[21] ;
 wire \wbd_mbist7_dat_o[22] ;
 wire \wbd_mbist7_dat_o[23] ;
 wire \wbd_mbist7_dat_o[24] ;
 wire \wbd_mbist7_dat_o[25] ;
 wire \wbd_mbist7_dat_o[26] ;
 wire \wbd_mbist7_dat_o[27] ;
 wire \wbd_mbist7_dat_o[28] ;
 wire \wbd_mbist7_dat_o[29] ;
 wire \wbd_mbist7_dat_o[2] ;
 wire \wbd_mbist7_dat_o[30] ;
 wire \wbd_mbist7_dat_o[31] ;
 wire \wbd_mbist7_dat_o[3] ;
 wire \wbd_mbist7_dat_o[4] ;
 wire \wbd_mbist7_dat_o[5] ;
 wire \wbd_mbist7_dat_o[6] ;
 wire \wbd_mbist7_dat_o[7] ;
 wire \wbd_mbist7_dat_o[8] ;
 wire \wbd_mbist7_dat_o[9] ;
 wire \wbd_mbist7_sel_o[0] ;
 wire \wbd_mbist7_sel_o[1] ;
 wire \wbd_mbist7_sel_o[2] ;
 wire \wbd_mbist7_sel_o[3] ;
 wire wbd_mbist7_stb_o;
 wire wbd_mbist7_we_o;
 wire wbd_mbist8_ack_i;
 wire \wbd_mbist8_adr_o[0] ;
 wire \wbd_mbist8_adr_o[1] ;
 wire \wbd_mbist8_adr_o[2] ;
 wire \wbd_mbist8_adr_o[3] ;
 wire \wbd_mbist8_adr_o[4] ;
 wire \wbd_mbist8_adr_o[5] ;
 wire \wbd_mbist8_adr_o[6] ;
 wire \wbd_mbist8_adr_o[7] ;
 wire \wbd_mbist8_adr_o[8] ;
 wire \wbd_mbist8_adr_o[9] ;
 wire wbd_mbist8_cyc_o;
 wire \wbd_mbist8_dat_i[0] ;
 wire \wbd_mbist8_dat_i[10] ;
 wire \wbd_mbist8_dat_i[11] ;
 wire \wbd_mbist8_dat_i[12] ;
 wire \wbd_mbist8_dat_i[13] ;
 wire \wbd_mbist8_dat_i[14] ;
 wire \wbd_mbist8_dat_i[15] ;
 wire \wbd_mbist8_dat_i[16] ;
 wire \wbd_mbist8_dat_i[17] ;
 wire \wbd_mbist8_dat_i[18] ;
 wire \wbd_mbist8_dat_i[19] ;
 wire \wbd_mbist8_dat_i[1] ;
 wire \wbd_mbist8_dat_i[20] ;
 wire \wbd_mbist8_dat_i[21] ;
 wire \wbd_mbist8_dat_i[22] ;
 wire \wbd_mbist8_dat_i[23] ;
 wire \wbd_mbist8_dat_i[24] ;
 wire \wbd_mbist8_dat_i[25] ;
 wire \wbd_mbist8_dat_i[26] ;
 wire \wbd_mbist8_dat_i[27] ;
 wire \wbd_mbist8_dat_i[28] ;
 wire \wbd_mbist8_dat_i[29] ;
 wire \wbd_mbist8_dat_i[2] ;
 wire \wbd_mbist8_dat_i[30] ;
 wire \wbd_mbist8_dat_i[31] ;
 wire \wbd_mbist8_dat_i[3] ;
 wire \wbd_mbist8_dat_i[4] ;
 wire \wbd_mbist8_dat_i[5] ;
 wire \wbd_mbist8_dat_i[6] ;
 wire \wbd_mbist8_dat_i[7] ;
 wire \wbd_mbist8_dat_i[8] ;
 wire \wbd_mbist8_dat_i[9] ;
 wire \wbd_mbist8_dat_o[0] ;
 wire \wbd_mbist8_dat_o[10] ;
 wire \wbd_mbist8_dat_o[11] ;
 wire \wbd_mbist8_dat_o[12] ;
 wire \wbd_mbist8_dat_o[13] ;
 wire \wbd_mbist8_dat_o[14] ;
 wire \wbd_mbist8_dat_o[15] ;
 wire \wbd_mbist8_dat_o[16] ;
 wire \wbd_mbist8_dat_o[17] ;
 wire \wbd_mbist8_dat_o[18] ;
 wire \wbd_mbist8_dat_o[19] ;
 wire \wbd_mbist8_dat_o[1] ;
 wire \wbd_mbist8_dat_o[20] ;
 wire \wbd_mbist8_dat_o[21] ;
 wire \wbd_mbist8_dat_o[22] ;
 wire \wbd_mbist8_dat_o[23] ;
 wire \wbd_mbist8_dat_o[24] ;
 wire \wbd_mbist8_dat_o[25] ;
 wire \wbd_mbist8_dat_o[26] ;
 wire \wbd_mbist8_dat_o[27] ;
 wire \wbd_mbist8_dat_o[28] ;
 wire \wbd_mbist8_dat_o[29] ;
 wire \wbd_mbist8_dat_o[2] ;
 wire \wbd_mbist8_dat_o[30] ;
 wire \wbd_mbist8_dat_o[31] ;
 wire \wbd_mbist8_dat_o[3] ;
 wire \wbd_mbist8_dat_o[4] ;
 wire \wbd_mbist8_dat_o[5] ;
 wire \wbd_mbist8_dat_o[6] ;
 wire \wbd_mbist8_dat_o[7] ;
 wire \wbd_mbist8_dat_o[8] ;
 wire \wbd_mbist8_dat_o[9] ;
 wire \wbd_mbist8_sel_o[0] ;
 wire \wbd_mbist8_sel_o[1] ;
 wire \wbd_mbist8_sel_o[2] ;
 wire \wbd_mbist8_sel_o[3] ;
 wire wbd_mbist8_stb_o;
 wire wbd_mbist8_we_o;

 glbl_cfg u_glbl (.mclk(wbd_clk_glbl),
    .reg_ack(wbd_glbl_ack_i),
    .reg_cs(wbd_glbl_stb_o),
    .reg_wr(wbd_glbl_we_o),
    .reset_n(wbd_int_rst_n),
    .scan_en(scan_en),
    .scan_en_o(scan_en_glbl),
    .scan_mode(scan_mode),
    .scan_mode_o(scan_mode_glbl),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbd_clk_glbl(wbd_clk_glbl),
    .wbd_clk_int(wbd_clk_glbl_int),
    .bist_correct({\bist_correct_int[7] ,
    \bist_correct_int[6] ,
    \bist_correct_int[5] ,
    \bist_correct_int[4] ,
    \bist_correct_int[3] ,
    \bist_correct_int[2] ,
    \bist_correct_int[1] ,
    \bist_correct_int[0] }),
    .bist_done({\bist_done_int[7] ,
    \bist_done_int[6] ,
    \bist_done_int[5] ,
    \bist_done_int[4] ,
    \bist_done_int[3] ,
    \bist_done_int[2] ,
    \bist_done_int[1] ,
    \bist_done_int[0] }),
    .bist_en({\bist_en[7] ,
    \bist_en[6] ,
    \bist_en[5] ,
    \bist_en[4] ,
    \bist_en[3] ,
    \bist_en[2] ,
    \bist_en[1] ,
    \bist_en[0] }),
    .bist_error({\bist_error_int[7] ,
    \bist_error_int[6] ,
    \bist_error_int[5] ,
    \bist_error_int[4] ,
    \bist_error_int[3] ,
    \bist_error_int[2] ,
    \bist_error_int[1] ,
    \bist_error_int[0] }),
    .bist_error_cnt0({\bist_error_cnt0_int[3] ,
    \bist_error_cnt0_int[2] ,
    \bist_error_cnt0_int[1] ,
    \bist_error_cnt0_int[0] }),
    .bist_error_cnt1({\bist_error_cnt1_int[3] ,
    \bist_error_cnt1_int[2] ,
    \bist_error_cnt1_int[1] ,
    \bist_error_cnt1_int[0] }),
    .bist_error_cnt2({\bist_error_cnt2_int[3] ,
    \bist_error_cnt2_int[2] ,
    \bist_error_cnt2_int[1] ,
    \bist_error_cnt2_int[0] }),
    .bist_error_cnt3({\bist_error_cnt3_int[3] ,
    \bist_error_cnt3_int[2] ,
    \bist_error_cnt3_int[1] ,
    \bist_error_cnt3_int[0] }),
    .bist_error_cnt4({\bist_error_cnt4_int[3] ,
    \bist_error_cnt4_int[2] ,
    \bist_error_cnt4_int[1] ,
    \bist_error_cnt4_int[0] }),
    .bist_error_cnt5({\bist_error_cnt5_int[3] ,
    \bist_error_cnt5_int[2] ,
    \bist_error_cnt5_int[1] ,
    \bist_error_cnt5_int[0] }),
    .bist_error_cnt6({\bist_error_cnt6_int[3] ,
    \bist_error_cnt6_int[2] ,
    \bist_error_cnt6_int[1] ,
    \bist_error_cnt6_int[0] }),
    .bist_error_cnt7({\bist_error_cnt7_int[3] ,
    \bist_error_cnt7_int[2] ,
    \bist_error_cnt7_int[1] ,
    \bist_error_cnt7_int[0] }),
    .bist_load({\bist_load[7] ,
    \bist_load[6] ,
    \bist_load[5] ,
    \bist_load[4] ,
    \bist_load[3] ,
    \bist_load[2] ,
    \bist_load[1] ,
    \bist_load[0] }),
    .bist_run({\bist_run[7] ,
    \bist_run[6] ,
    \bist_run[5] ,
    \bist_run[4] ,
    \bist_run[3] ,
    \bist_run[2] ,
    \bist_run[1] ,
    \bist_run[0] }),
    .bist_sdi({\bist_sdi[7] ,
    \bist_sdi[6] ,
    \bist_sdi[5] ,
    \bist_sdi[4] ,
    \bist_sdi[3] ,
    \bist_sdi[2] ,
    \bist_sdi[1] ,
    \bist_sdi[0] }),
    .bist_sdo({\bist_sdo_int[7] ,
    \bist_sdo_int[6] ,
    \bist_sdo_int[5] ,
    \bist_sdo_int[4] ,
    \bist_sdo_int[3] ,
    \bist_sdo_int[2] ,
    \bist_sdo_int[1] ,
    \bist_sdo_int[0] }),
    .bist_shift({\bist_shift[7] ,
    \bist_shift[6] ,
    \bist_shift[5] ,
    \bist_shift[4] ,
    \bist_shift[3] ,
    \bist_shift[2] ,
    \bist_shift[1] ,
    \bist_shift[0] }),
    .cfg_cska_glbl({\cfg_clk_ctrl1[11] ,
    \cfg_clk_ctrl1[10] ,
    \cfg_clk_ctrl1[9] ,
    \cfg_clk_ctrl1[8] }),
    .reg_addr({\wbd_glbl_adr_o[7] ,
    \wbd_glbl_adr_o[6] ,
    \wbd_glbl_adr_o[5] ,
    \wbd_glbl_adr_o[4] ,
    \wbd_glbl_adr_o[3] ,
    \wbd_glbl_adr_o[2] ,
    \wbd_glbl_adr_o[1] ,
    \wbd_glbl_adr_o[0] }),
    .reg_be({\wbd_glbl_sel_o[3] ,
    \wbd_glbl_sel_o[2] ,
    \wbd_glbl_sel_o[1] ,
    \wbd_glbl_sel_o[0] }),
    .reg_rdata({\wbd_glbl_dat_i[31] ,
    \wbd_glbl_dat_i[30] ,
    \wbd_glbl_dat_i[29] ,
    \wbd_glbl_dat_i[28] ,
    \wbd_glbl_dat_i[27] ,
    \wbd_glbl_dat_i[26] ,
    \wbd_glbl_dat_i[25] ,
    \wbd_glbl_dat_i[24] ,
    \wbd_glbl_dat_i[23] ,
    \wbd_glbl_dat_i[22] ,
    \wbd_glbl_dat_i[21] ,
    \wbd_glbl_dat_i[20] ,
    \wbd_glbl_dat_i[19] ,
    \wbd_glbl_dat_i[18] ,
    \wbd_glbl_dat_i[17] ,
    \wbd_glbl_dat_i[16] ,
    \wbd_glbl_dat_i[15] ,
    \wbd_glbl_dat_i[14] ,
    \wbd_glbl_dat_i[13] ,
    \wbd_glbl_dat_i[12] ,
    \wbd_glbl_dat_i[11] ,
    \wbd_glbl_dat_i[10] ,
    \wbd_glbl_dat_i[9] ,
    \wbd_glbl_dat_i[8] ,
    \wbd_glbl_dat_i[7] ,
    \wbd_glbl_dat_i[6] ,
    \wbd_glbl_dat_i[5] ,
    \wbd_glbl_dat_i[4] ,
    \wbd_glbl_dat_i[3] ,
    \wbd_glbl_dat_i[2] ,
    \wbd_glbl_dat_i[1] ,
    \wbd_glbl_dat_i[0] }),
    .reg_wdata({\wbd_glbl_dat_o[31] ,
    \wbd_glbl_dat_o[30] ,
    \wbd_glbl_dat_o[29] ,
    \wbd_glbl_dat_o[28] ,
    \wbd_glbl_dat_o[27] ,
    \wbd_glbl_dat_o[26] ,
    \wbd_glbl_dat_o[25] ,
    \wbd_glbl_dat_o[24] ,
    \wbd_glbl_dat_o[23] ,
    \wbd_glbl_dat_o[22] ,
    \wbd_glbl_dat_o[21] ,
    \wbd_glbl_dat_o[20] ,
    \wbd_glbl_dat_o[19] ,
    \wbd_glbl_dat_o[18] ,
    \wbd_glbl_dat_o[17] ,
    \wbd_glbl_dat_o[16] ,
    \wbd_glbl_dat_o[15] ,
    \wbd_glbl_dat_o[14] ,
    \wbd_glbl_dat_o[13] ,
    \wbd_glbl_dat_o[12] ,
    \wbd_glbl_dat_o[11] ,
    \wbd_glbl_dat_o[10] ,
    \wbd_glbl_dat_o[9] ,
    \wbd_glbl_dat_o[8] ,
    \wbd_glbl_dat_o[7] ,
    \wbd_glbl_dat_o[6] ,
    \wbd_glbl_dat_o[5] ,
    \wbd_glbl_dat_o[4] ,
    \wbd_glbl_dat_o[3] ,
    \wbd_glbl_dat_o[2] ,
    \wbd_glbl_dat_o[1] ,
    \wbd_glbl_dat_o[0] }),
    .scan_si({\scan_in[7] ,
    \scan_in[6] ,
    \scan_in[5] ,
    \scan_in[4] ,
    \scan_in[3] ,
    \scan_in[2] ,
    \scan_in[1] ,
    \scan_in[0] }),
    .scan_so({\scan_out_glbl[7] ,
    \scan_out_glbl[6] ,
    \scan_out_glbl[5] ,
    \scan_out_glbl[4] ,
    \scan_out_glbl[3] ,
    \scan_out_glbl[2] ,
    \scan_out_glbl[1] ,
    \scan_out_glbl[0] }));
 wb_interconnect u_intercon (.clk_i(wbd_clk_wi),
    .m0_wbd_ack_o(wbd_int_ack_o),
    .m0_wbd_cyc_i(wbd_int_cyc_i),
    .m0_wbd_err_o(wbd_int_err_o),
    .m0_wbd_stb_i(wbd_int_stb_i),
    .m0_wbd_we_i(wbd_int_we_i),
    .rst_n(wbd_int_rst_n),
    .s0_wbd_ack_i(wbd_glbl_ack_i),
    .s0_wbd_cyc_o(wbd_glbl_cyc_o),
    .s0_wbd_stb_o(wbd_glbl_stb_o),
    .s0_wbd_we_o(wbd_glbl_we_o),
    .s1_wbd_ack_i(wbd_mbist1_ack_i),
    .s1_wbd_cyc_o(wbd_mbist1_cyc_o),
    .s1_wbd_stb_o(wbd_mbist1_stb_o),
    .s1_wbd_we_o(wbd_mbist1_we_o),
    .s2_wbd_ack_i(wbd_mbist2_ack_i),
    .s2_wbd_cyc_o(wbd_mbist2_cyc_o),
    .s2_wbd_stb_o(wbd_mbist2_stb_o),
    .s2_wbd_we_o(wbd_mbist2_we_o),
    .s3_wbd_ack_i(wbd_mbist3_ack_i),
    .s3_wbd_cyc_o(wbd_mbist3_cyc_o),
    .s3_wbd_stb_o(wbd_mbist3_stb_o),
    .s3_wbd_we_o(wbd_mbist3_we_o),
    .s4_wbd_ack_i(wbd_mbist4_ack_i),
    .s4_wbd_cyc_o(wbd_mbist4_cyc_o),
    .s4_wbd_stb_o(wbd_mbist4_stb_o),
    .s4_wbd_we_o(wbd_mbist4_we_o),
    .s5_wbd_ack_i(wbd_mbist5_ack_i),
    .s5_wbd_cyc_o(wbd_mbist5_cyc_o),
    .s5_wbd_stb_o(wbd_mbist5_stb_o),
    .s5_wbd_we_o(wbd_mbist5_we_o),
    .s6_wbd_ack_i(wbd_mbist6_ack_i),
    .s6_wbd_cyc_o(wbd_mbist6_cyc_o),
    .s6_wbd_stb_o(wbd_mbist6_stb_o),
    .s6_wbd_we_o(wbd_mbist6_we_o),
    .s7_wbd_ack_i(wbd_mbist7_ack_i),
    .s7_wbd_cyc_o(wbd_mbist7_cyc_o),
    .s7_wbd_stb_o(wbd_mbist7_stb_o),
    .s7_wbd_we_o(wbd_mbist7_we_o),
    .s8_wbd_ack_i(wbd_mbist8_ack_i),
    .s8_wbd_cyc_o(wbd_mbist8_cyc_o),
    .s8_wbd_stb_o(wbd_mbist8_stb_o),
    .s8_wbd_we_o(wbd_mbist8_we_o),
    .scan_en(scan_en_mbist8),
    .scan_en_o(scan_en_wbi),
    .scan_mode(scan_mode_mbist8),
    .scan_mode_o(scan_mode_wbi),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbd_clk_int(wbd_clk_int),
    .wbd_clk_wi(wbd_clk_wi),
    .cfg_cska_wi({\cfg_clk_ctrl1[7] ,
    \cfg_clk_ctrl1[6] ,
    \cfg_clk_ctrl1[5] ,
    \cfg_clk_ctrl1[4] }),
    .ch_clk_in({wbd_clk_int,
    wbd_clk_int,
    wbd_clk_int,
    wbd_clk_int,
    wbd_clk_int,
    wbd_clk_int,
    wbd_clk_int,
    wbd_clk_int,
    wbd_clk_int}),
    .ch_clk_out({wbd_clk_mbist8_int,
    wbd_clk_mbist7_int,
    wbd_clk_mbist6_int,
    wbd_clk_mbist5_int,
    wbd_clk_mbist4_int,
    wbd_clk_mbist3_int,
    wbd_clk_mbist2_int,
    wbd_clk_mbist1_int,
    wbd_clk_glbl_int}),
    .ch_data_in({\bist_error_cnt7[3] ,
    \bist_error_cnt7[2] ,
    \bist_error_cnt7[1] ,
    \bist_error_cnt7[0] ,
    \bist_correct[7] ,
    \bist_error[7] ,
    \bist_done[7] ,
    \bist_sdo[7] ,
    \bist_sdi[7] ,
    \bist_load[7] ,
    \bist_shift[7] ,
    \bist_run[7] ,
    \bist_en[7] ,
    \bist_error_cnt6[3] ,
    \bist_error_cnt6[2] ,
    \bist_error_cnt6[1] ,
    \bist_error_cnt6[0] ,
    \bist_correct[6] ,
    \bist_error[6] ,
    \bist_done[6] ,
    \bist_sdo[6] ,
    \bist_sdi[6] ,
    \bist_load[6] ,
    \bist_shift[6] ,
    \bist_run[6] ,
    \bist_en[6] ,
    \bist_error_cnt5[3] ,
    \bist_error_cnt5[2] ,
    \bist_error_cnt5[1] ,
    \bist_error_cnt5[0] ,
    \bist_correct[5] ,
    \bist_error[5] ,
    \bist_done[5] ,
    \bist_sdo[5] ,
    \bist_sdi[5] ,
    \bist_load[5] ,
    \bist_shift[5] ,
    \bist_run[5] ,
    \bist_en[5] ,
    \bist_error_cnt4[3] ,
    \bist_error_cnt4[2] ,
    \bist_error_cnt4[1] ,
    \bist_error_cnt4[0] ,
    \bist_correct[4] ,
    \bist_error[4] ,
    \bist_done[4] ,
    \bist_sdo[4] ,
    \bist_sdi[4] ,
    \bist_load[4] ,
    \bist_shift[4] ,
    \bist_run[4] ,
    \bist_en[4] ,
    \bist_error_cnt3[3] ,
    \bist_error_cnt3[2] ,
    \bist_error_cnt3[1] ,
    \bist_error_cnt3[0] ,
    \bist_correct[3] ,
    \bist_error[3] ,
    \bist_done[3] ,
    \bist_sdo[3] ,
    \bist_sdi[3] ,
    \bist_load[3] ,
    \bist_shift[3] ,
    \bist_run[3] ,
    \bist_en[3] ,
    \bist_error_cnt2[3] ,
    \bist_error_cnt2[2] ,
    \bist_error_cnt2[1] ,
    \bist_error_cnt2[0] ,
    \bist_correct[2] ,
    \bist_error[2] ,
    \bist_done[2] ,
    \bist_sdo[2] ,
    \bist_sdi[2] ,
    \bist_load[2] ,
    \bist_shift[2] ,
    \bist_run[2] ,
    \bist_en[2] ,
    \bist_error_cnt1[3] ,
    \bist_error_cnt1[2] ,
    \bist_error_cnt1[1] ,
    \bist_error_cnt1[0] ,
    \bist_correct[1] ,
    \bist_error[1] ,
    \bist_done[1] ,
    \bist_sdo[1] ,
    \bist_sdi[1] ,
    \bist_load[1] ,
    \bist_shift[1] ,
    \bist_run[1] ,
    \bist_en[1] ,
    \bist_error_cnt0[3] ,
    \bist_error_cnt0[2] ,
    \bist_error_cnt0[1] ,
    \bist_error_cnt0[0] ,
    \bist_correct[0] ,
    \bist_error[0] ,
    \bist_done[0] ,
    \bist_sdo[0] ,
    \bist_sdi[0] ,
    \bist_load[0] ,
    \bist_shift[0] ,
    \bist_run[0] ,
    \bist_en[0] }),
    .ch_data_out({\bist_error_cnt7_int[3] ,
    \bist_error_cnt7_int[2] ,
    \bist_error_cnt7_int[1] ,
    \bist_error_cnt7_int[0] ,
    \bist_correct_int[7] ,
    \bist_error_int[7] ,
    \bist_done_int[7] ,
    \bist_sdo_int[7] ,
    \bist_sdi_int[7] ,
    \bist_load_int[7] ,
    \bist_shift_int[7] ,
    \bist_run_int[7] ,
    \bist_en_int[7] ,
    \bist_error_cnt6_int[3] ,
    \bist_error_cnt6_int[2] ,
    \bist_error_cnt6_int[1] ,
    \bist_error_cnt6_int[0] ,
    \bist_correct_int[6] ,
    \bist_error_int[6] ,
    \bist_done_int[6] ,
    \bist_sdo_int[6] ,
    \bist_sdi_int[6] ,
    \bist_load_int[6] ,
    \bist_shift_int[6] ,
    \bist_run_int[6] ,
    \bist_en_int[6] ,
    \bist_error_cnt5_int[3] ,
    \bist_error_cnt5_int[2] ,
    \bist_error_cnt5_int[1] ,
    \bist_error_cnt5_int[0] ,
    \bist_correct_int[5] ,
    \bist_error_int[5] ,
    \bist_done_int[5] ,
    \bist_sdo_int[5] ,
    \bist_sdi_int[5] ,
    \bist_load_int[5] ,
    \bist_shift_int[5] ,
    \bist_run_int[5] ,
    \bist_en_int[5] ,
    \bist_error_cnt4_int[3] ,
    \bist_error_cnt4_int[2] ,
    \bist_error_cnt4_int[1] ,
    \bist_error_cnt4_int[0] ,
    \bist_correct_int[4] ,
    \bist_error_int[4] ,
    \bist_done_int[4] ,
    \bist_sdo_int[4] ,
    \bist_sdi_int[4] ,
    \bist_load_int[4] ,
    \bist_shift_int[4] ,
    \bist_run_int[4] ,
    \bist_en_int[4] ,
    \bist_error_cnt3_int[3] ,
    \bist_error_cnt3_int[2] ,
    \bist_error_cnt3_int[1] ,
    \bist_error_cnt3_int[0] ,
    \bist_correct_int[3] ,
    \bist_error_int[3] ,
    \bist_done_int[3] ,
    \bist_sdo_int[3] ,
    \bist_sdi_int[3] ,
    \bist_load_int[3] ,
    \bist_shift_int[3] ,
    \bist_run_int[3] ,
    \bist_en_int[3] ,
    \bist_error_cnt2_int[3] ,
    \bist_error_cnt2_int[2] ,
    \bist_error_cnt2_int[1] ,
    \bist_error_cnt2_int[0] ,
    \bist_correct_int[2] ,
    \bist_error_int[2] ,
    \bist_done_int[2] ,
    \bist_sdo_int[2] ,
    \bist_sdi_int[2] ,
    \bist_load_int[2] ,
    \bist_shift_int[2] ,
    \bist_run_int[2] ,
    \bist_en_int[2] ,
    \bist_error_cnt1_int[3] ,
    \bist_error_cnt1_int[2] ,
    \bist_error_cnt1_int[1] ,
    \bist_error_cnt1_int[0] ,
    \bist_correct_int[1] ,
    \bist_error_int[1] ,
    \bist_done_int[1] ,
    \bist_sdo_int[1] ,
    \bist_sdi_int[1] ,
    \bist_load_int[1] ,
    \bist_shift_int[1] ,
    \bist_run_int[1] ,
    \bist_en_int[1] ,
    \bist_error_cnt0_int[3] ,
    \bist_error_cnt0_int[2] ,
    \bist_error_cnt0_int[1] ,
    \bist_error_cnt0_int[0] ,
    \bist_correct_int[0] ,
    \bist_error_int[0] ,
    \bist_done_int[0] ,
    \bist_sdo_int[0] ,
    \bist_sdi_int[0] ,
    \bist_load_int[0] ,
    \bist_shift_int[0] ,
    \bist_run_int[0] ,
    \bist_en_int[0] }),
    .m0_wbd_adr_i({\wbd_int_adr_i[31] ,
    \wbd_int_adr_i[30] ,
    \wbd_int_adr_i[29] ,
    \wbd_int_adr_i[28] ,
    \wbd_int_adr_i[27] ,
    \wbd_int_adr_i[26] ,
    \wbd_int_adr_i[25] ,
    \wbd_int_adr_i[24] ,
    \wbd_int_adr_i[23] ,
    \wbd_int_adr_i[22] ,
    \wbd_int_adr_i[21] ,
    \wbd_int_adr_i[20] ,
    \wbd_int_adr_i[19] ,
    \wbd_int_adr_i[18] ,
    \wbd_int_adr_i[17] ,
    \wbd_int_adr_i[16] ,
    \wbd_int_adr_i[15] ,
    \wbd_int_adr_i[14] ,
    \wbd_int_adr_i[13] ,
    \wbd_int_adr_i[12] ,
    \wbd_int_adr_i[11] ,
    \wbd_int_adr_i[10] ,
    \wbd_int_adr_i[9] ,
    \wbd_int_adr_i[8] ,
    \wbd_int_adr_i[7] ,
    \wbd_int_adr_i[6] ,
    \wbd_int_adr_i[5] ,
    \wbd_int_adr_i[4] ,
    \wbd_int_adr_i[3] ,
    \wbd_int_adr_i[2] ,
    \wbd_int_adr_i[1] ,
    \wbd_int_adr_i[0] }),
    .m0_wbd_dat_i({\wbd_int_dat_i[31] ,
    \wbd_int_dat_i[30] ,
    \wbd_int_dat_i[29] ,
    \wbd_int_dat_i[28] ,
    \wbd_int_dat_i[27] ,
    \wbd_int_dat_i[26] ,
    \wbd_int_dat_i[25] ,
    \wbd_int_dat_i[24] ,
    \wbd_int_dat_i[23] ,
    \wbd_int_dat_i[22] ,
    \wbd_int_dat_i[21] ,
    \wbd_int_dat_i[20] ,
    \wbd_int_dat_i[19] ,
    \wbd_int_dat_i[18] ,
    \wbd_int_dat_i[17] ,
    \wbd_int_dat_i[16] ,
    \wbd_int_dat_i[15] ,
    \wbd_int_dat_i[14] ,
    \wbd_int_dat_i[13] ,
    \wbd_int_dat_i[12] ,
    \wbd_int_dat_i[11] ,
    \wbd_int_dat_i[10] ,
    \wbd_int_dat_i[9] ,
    \wbd_int_dat_i[8] ,
    \wbd_int_dat_i[7] ,
    \wbd_int_dat_i[6] ,
    \wbd_int_dat_i[5] ,
    \wbd_int_dat_i[4] ,
    \wbd_int_dat_i[3] ,
    \wbd_int_dat_i[2] ,
    \wbd_int_dat_i[1] ,
    \wbd_int_dat_i[0] }),
    .m0_wbd_dat_o({\wbd_int_dat_o[31] ,
    \wbd_int_dat_o[30] ,
    \wbd_int_dat_o[29] ,
    \wbd_int_dat_o[28] ,
    \wbd_int_dat_o[27] ,
    \wbd_int_dat_o[26] ,
    \wbd_int_dat_o[25] ,
    \wbd_int_dat_o[24] ,
    \wbd_int_dat_o[23] ,
    \wbd_int_dat_o[22] ,
    \wbd_int_dat_o[21] ,
    \wbd_int_dat_o[20] ,
    \wbd_int_dat_o[19] ,
    \wbd_int_dat_o[18] ,
    \wbd_int_dat_o[17] ,
    \wbd_int_dat_o[16] ,
    \wbd_int_dat_o[15] ,
    \wbd_int_dat_o[14] ,
    \wbd_int_dat_o[13] ,
    \wbd_int_dat_o[12] ,
    \wbd_int_dat_o[11] ,
    \wbd_int_dat_o[10] ,
    \wbd_int_dat_o[9] ,
    \wbd_int_dat_o[8] ,
    \wbd_int_dat_o[7] ,
    \wbd_int_dat_o[6] ,
    \wbd_int_dat_o[5] ,
    \wbd_int_dat_o[4] ,
    \wbd_int_dat_o[3] ,
    \wbd_int_dat_o[2] ,
    \wbd_int_dat_o[1] ,
    \wbd_int_dat_o[0] }),
    .m0_wbd_sel_i({\wbd_int_sel_i[3] ,
    \wbd_int_sel_i[2] ,
    \wbd_int_sel_i[1] ,
    \wbd_int_sel_i[0] }),
    .s0_wbd_adr_o({\wbd_glbl_adr_o[7] ,
    \wbd_glbl_adr_o[6] ,
    \wbd_glbl_adr_o[5] ,
    \wbd_glbl_adr_o[4] ,
    \wbd_glbl_adr_o[3] ,
    \wbd_glbl_adr_o[2] ,
    \wbd_glbl_adr_o[1] ,
    \wbd_glbl_adr_o[0] }),
    .s0_wbd_dat_i({\wbd_glbl_dat_i[31] ,
    \wbd_glbl_dat_i[30] ,
    \wbd_glbl_dat_i[29] ,
    \wbd_glbl_dat_i[28] ,
    \wbd_glbl_dat_i[27] ,
    \wbd_glbl_dat_i[26] ,
    \wbd_glbl_dat_i[25] ,
    \wbd_glbl_dat_i[24] ,
    \wbd_glbl_dat_i[23] ,
    \wbd_glbl_dat_i[22] ,
    \wbd_glbl_dat_i[21] ,
    \wbd_glbl_dat_i[20] ,
    \wbd_glbl_dat_i[19] ,
    \wbd_glbl_dat_i[18] ,
    \wbd_glbl_dat_i[17] ,
    \wbd_glbl_dat_i[16] ,
    \wbd_glbl_dat_i[15] ,
    \wbd_glbl_dat_i[14] ,
    \wbd_glbl_dat_i[13] ,
    \wbd_glbl_dat_i[12] ,
    \wbd_glbl_dat_i[11] ,
    \wbd_glbl_dat_i[10] ,
    \wbd_glbl_dat_i[9] ,
    \wbd_glbl_dat_i[8] ,
    \wbd_glbl_dat_i[7] ,
    \wbd_glbl_dat_i[6] ,
    \wbd_glbl_dat_i[5] ,
    \wbd_glbl_dat_i[4] ,
    \wbd_glbl_dat_i[3] ,
    \wbd_glbl_dat_i[2] ,
    \wbd_glbl_dat_i[1] ,
    \wbd_glbl_dat_i[0] }),
    .s0_wbd_dat_o({\wbd_glbl_dat_o[31] ,
    \wbd_glbl_dat_o[30] ,
    \wbd_glbl_dat_o[29] ,
    \wbd_glbl_dat_o[28] ,
    \wbd_glbl_dat_o[27] ,
    \wbd_glbl_dat_o[26] ,
    \wbd_glbl_dat_o[25] ,
    \wbd_glbl_dat_o[24] ,
    \wbd_glbl_dat_o[23] ,
    \wbd_glbl_dat_o[22] ,
    \wbd_glbl_dat_o[21] ,
    \wbd_glbl_dat_o[20] ,
    \wbd_glbl_dat_o[19] ,
    \wbd_glbl_dat_o[18] ,
    \wbd_glbl_dat_o[17] ,
    \wbd_glbl_dat_o[16] ,
    \wbd_glbl_dat_o[15] ,
    \wbd_glbl_dat_o[14] ,
    \wbd_glbl_dat_o[13] ,
    \wbd_glbl_dat_o[12] ,
    \wbd_glbl_dat_o[11] ,
    \wbd_glbl_dat_o[10] ,
    \wbd_glbl_dat_o[9] ,
    \wbd_glbl_dat_o[8] ,
    \wbd_glbl_dat_o[7] ,
    \wbd_glbl_dat_o[6] ,
    \wbd_glbl_dat_o[5] ,
    \wbd_glbl_dat_o[4] ,
    \wbd_glbl_dat_o[3] ,
    \wbd_glbl_dat_o[2] ,
    \wbd_glbl_dat_o[1] ,
    \wbd_glbl_dat_o[0] }),
    .s0_wbd_sel_o({\wbd_glbl_sel_o[3] ,
    \wbd_glbl_sel_o[2] ,
    \wbd_glbl_sel_o[1] ,
    \wbd_glbl_sel_o[0] }),
    .s1_wbd_adr_o({\wbd_mbist1_adr_o[10] ,
    \wbd_mbist1_adr_o[9] ,
    \wbd_mbist1_adr_o[8] ,
    \wbd_mbist1_adr_o[7] ,
    \wbd_mbist1_adr_o[6] ,
    \wbd_mbist1_adr_o[5] ,
    \wbd_mbist1_adr_o[4] ,
    \wbd_mbist1_adr_o[3] ,
    \wbd_mbist1_adr_o[2] ,
    \wbd_mbist1_adr_o[1] ,
    \wbd_mbist1_adr_o[0] }),
    .s1_wbd_dat_i({\wbd_mbist1_dat_i[31] ,
    \wbd_mbist1_dat_i[30] ,
    \wbd_mbist1_dat_i[29] ,
    \wbd_mbist1_dat_i[28] ,
    \wbd_mbist1_dat_i[27] ,
    \wbd_mbist1_dat_i[26] ,
    \wbd_mbist1_dat_i[25] ,
    \wbd_mbist1_dat_i[24] ,
    \wbd_mbist1_dat_i[23] ,
    \wbd_mbist1_dat_i[22] ,
    \wbd_mbist1_dat_i[21] ,
    \wbd_mbist1_dat_i[20] ,
    \wbd_mbist1_dat_i[19] ,
    \wbd_mbist1_dat_i[18] ,
    \wbd_mbist1_dat_i[17] ,
    \wbd_mbist1_dat_i[16] ,
    \wbd_mbist1_dat_i[15] ,
    \wbd_mbist1_dat_i[14] ,
    \wbd_mbist1_dat_i[13] ,
    \wbd_mbist1_dat_i[12] ,
    \wbd_mbist1_dat_i[11] ,
    \wbd_mbist1_dat_i[10] ,
    \wbd_mbist1_dat_i[9] ,
    \wbd_mbist1_dat_i[8] ,
    \wbd_mbist1_dat_i[7] ,
    \wbd_mbist1_dat_i[6] ,
    \wbd_mbist1_dat_i[5] ,
    \wbd_mbist1_dat_i[4] ,
    \wbd_mbist1_dat_i[3] ,
    \wbd_mbist1_dat_i[2] ,
    \wbd_mbist1_dat_i[1] ,
    \wbd_mbist1_dat_i[0] }),
    .s1_wbd_dat_o({\wbd_mbist1_dat_o[31] ,
    \wbd_mbist1_dat_o[30] ,
    \wbd_mbist1_dat_o[29] ,
    \wbd_mbist1_dat_o[28] ,
    \wbd_mbist1_dat_o[27] ,
    \wbd_mbist1_dat_o[26] ,
    \wbd_mbist1_dat_o[25] ,
    \wbd_mbist1_dat_o[24] ,
    \wbd_mbist1_dat_o[23] ,
    \wbd_mbist1_dat_o[22] ,
    \wbd_mbist1_dat_o[21] ,
    \wbd_mbist1_dat_o[20] ,
    \wbd_mbist1_dat_o[19] ,
    \wbd_mbist1_dat_o[18] ,
    \wbd_mbist1_dat_o[17] ,
    \wbd_mbist1_dat_o[16] ,
    \wbd_mbist1_dat_o[15] ,
    \wbd_mbist1_dat_o[14] ,
    \wbd_mbist1_dat_o[13] ,
    \wbd_mbist1_dat_o[12] ,
    \wbd_mbist1_dat_o[11] ,
    \wbd_mbist1_dat_o[10] ,
    \wbd_mbist1_dat_o[9] ,
    \wbd_mbist1_dat_o[8] ,
    \wbd_mbist1_dat_o[7] ,
    \wbd_mbist1_dat_o[6] ,
    \wbd_mbist1_dat_o[5] ,
    \wbd_mbist1_dat_o[4] ,
    \wbd_mbist1_dat_o[3] ,
    \wbd_mbist1_dat_o[2] ,
    \wbd_mbist1_dat_o[1] ,
    \wbd_mbist1_dat_o[0] }),
    .s1_wbd_sel_o({\wbd_mbist1_sel_o[3] ,
    \wbd_mbist1_sel_o[2] ,
    \wbd_mbist1_sel_o[1] ,
    \wbd_mbist1_sel_o[0] }),
    .s2_wbd_adr_o({\wbd_mbist2_adr_o[10] ,
    \wbd_mbist2_adr_o[9] ,
    \wbd_mbist2_adr_o[8] ,
    \wbd_mbist2_adr_o[7] ,
    \wbd_mbist2_adr_o[6] ,
    \wbd_mbist2_adr_o[5] ,
    \wbd_mbist2_adr_o[4] ,
    \wbd_mbist2_adr_o[3] ,
    \wbd_mbist2_adr_o[2] ,
    \wbd_mbist2_adr_o[1] ,
    \wbd_mbist2_adr_o[0] }),
    .s2_wbd_dat_i({\wbd_mbist2_dat_i[31] ,
    \wbd_mbist2_dat_i[30] ,
    \wbd_mbist2_dat_i[29] ,
    \wbd_mbist2_dat_i[28] ,
    \wbd_mbist2_dat_i[27] ,
    \wbd_mbist2_dat_i[26] ,
    \wbd_mbist2_dat_i[25] ,
    \wbd_mbist2_dat_i[24] ,
    \wbd_mbist2_dat_i[23] ,
    \wbd_mbist2_dat_i[22] ,
    \wbd_mbist2_dat_i[21] ,
    \wbd_mbist2_dat_i[20] ,
    \wbd_mbist2_dat_i[19] ,
    \wbd_mbist2_dat_i[18] ,
    \wbd_mbist2_dat_i[17] ,
    \wbd_mbist2_dat_i[16] ,
    \wbd_mbist2_dat_i[15] ,
    \wbd_mbist2_dat_i[14] ,
    \wbd_mbist2_dat_i[13] ,
    \wbd_mbist2_dat_i[12] ,
    \wbd_mbist2_dat_i[11] ,
    \wbd_mbist2_dat_i[10] ,
    \wbd_mbist2_dat_i[9] ,
    \wbd_mbist2_dat_i[8] ,
    \wbd_mbist2_dat_i[7] ,
    \wbd_mbist2_dat_i[6] ,
    \wbd_mbist2_dat_i[5] ,
    \wbd_mbist2_dat_i[4] ,
    \wbd_mbist2_dat_i[3] ,
    \wbd_mbist2_dat_i[2] ,
    \wbd_mbist2_dat_i[1] ,
    \wbd_mbist2_dat_i[0] }),
    .s2_wbd_dat_o({\wbd_mbist2_dat_o[31] ,
    \wbd_mbist2_dat_o[30] ,
    \wbd_mbist2_dat_o[29] ,
    \wbd_mbist2_dat_o[28] ,
    \wbd_mbist2_dat_o[27] ,
    \wbd_mbist2_dat_o[26] ,
    \wbd_mbist2_dat_o[25] ,
    \wbd_mbist2_dat_o[24] ,
    \wbd_mbist2_dat_o[23] ,
    \wbd_mbist2_dat_o[22] ,
    \wbd_mbist2_dat_o[21] ,
    \wbd_mbist2_dat_o[20] ,
    \wbd_mbist2_dat_o[19] ,
    \wbd_mbist2_dat_o[18] ,
    \wbd_mbist2_dat_o[17] ,
    \wbd_mbist2_dat_o[16] ,
    \wbd_mbist2_dat_o[15] ,
    \wbd_mbist2_dat_o[14] ,
    \wbd_mbist2_dat_o[13] ,
    \wbd_mbist2_dat_o[12] ,
    \wbd_mbist2_dat_o[11] ,
    \wbd_mbist2_dat_o[10] ,
    \wbd_mbist2_dat_o[9] ,
    \wbd_mbist2_dat_o[8] ,
    \wbd_mbist2_dat_o[7] ,
    \wbd_mbist2_dat_o[6] ,
    \wbd_mbist2_dat_o[5] ,
    \wbd_mbist2_dat_o[4] ,
    \wbd_mbist2_dat_o[3] ,
    \wbd_mbist2_dat_o[2] ,
    \wbd_mbist2_dat_o[1] ,
    \wbd_mbist2_dat_o[0] }),
    .s2_wbd_sel_o({\wbd_mbist2_sel_o[3] ,
    \wbd_mbist2_sel_o[2] ,
    \wbd_mbist2_sel_o[1] ,
    \wbd_mbist2_sel_o[0] }),
    .s3_wbd_adr_o({\wbd_mbist3_adr_o[10] ,
    \wbd_mbist3_adr_o[9] ,
    \wbd_mbist3_adr_o[8] ,
    \wbd_mbist3_adr_o[7] ,
    \wbd_mbist3_adr_o[6] ,
    \wbd_mbist3_adr_o[5] ,
    \wbd_mbist3_adr_o[4] ,
    \wbd_mbist3_adr_o[3] ,
    \wbd_mbist3_adr_o[2] ,
    \wbd_mbist3_adr_o[1] ,
    \wbd_mbist3_adr_o[0] }),
    .s3_wbd_dat_i({\wbd_mbist3_dat_i[31] ,
    \wbd_mbist3_dat_i[30] ,
    \wbd_mbist3_dat_i[29] ,
    \wbd_mbist3_dat_i[28] ,
    \wbd_mbist3_dat_i[27] ,
    \wbd_mbist3_dat_i[26] ,
    \wbd_mbist3_dat_i[25] ,
    \wbd_mbist3_dat_i[24] ,
    \wbd_mbist3_dat_i[23] ,
    \wbd_mbist3_dat_i[22] ,
    \wbd_mbist3_dat_i[21] ,
    \wbd_mbist3_dat_i[20] ,
    \wbd_mbist3_dat_i[19] ,
    \wbd_mbist3_dat_i[18] ,
    \wbd_mbist3_dat_i[17] ,
    \wbd_mbist3_dat_i[16] ,
    \wbd_mbist3_dat_i[15] ,
    \wbd_mbist3_dat_i[14] ,
    \wbd_mbist3_dat_i[13] ,
    \wbd_mbist3_dat_i[12] ,
    \wbd_mbist3_dat_i[11] ,
    \wbd_mbist3_dat_i[10] ,
    \wbd_mbist3_dat_i[9] ,
    \wbd_mbist3_dat_i[8] ,
    \wbd_mbist3_dat_i[7] ,
    \wbd_mbist3_dat_i[6] ,
    \wbd_mbist3_dat_i[5] ,
    \wbd_mbist3_dat_i[4] ,
    \wbd_mbist3_dat_i[3] ,
    \wbd_mbist3_dat_i[2] ,
    \wbd_mbist3_dat_i[1] ,
    \wbd_mbist3_dat_i[0] }),
    .s3_wbd_dat_o({\wbd_mbist3_dat_o[31] ,
    \wbd_mbist3_dat_o[30] ,
    \wbd_mbist3_dat_o[29] ,
    \wbd_mbist3_dat_o[28] ,
    \wbd_mbist3_dat_o[27] ,
    \wbd_mbist3_dat_o[26] ,
    \wbd_mbist3_dat_o[25] ,
    \wbd_mbist3_dat_o[24] ,
    \wbd_mbist3_dat_o[23] ,
    \wbd_mbist3_dat_o[22] ,
    \wbd_mbist3_dat_o[21] ,
    \wbd_mbist3_dat_o[20] ,
    \wbd_mbist3_dat_o[19] ,
    \wbd_mbist3_dat_o[18] ,
    \wbd_mbist3_dat_o[17] ,
    \wbd_mbist3_dat_o[16] ,
    \wbd_mbist3_dat_o[15] ,
    \wbd_mbist3_dat_o[14] ,
    \wbd_mbist3_dat_o[13] ,
    \wbd_mbist3_dat_o[12] ,
    \wbd_mbist3_dat_o[11] ,
    \wbd_mbist3_dat_o[10] ,
    \wbd_mbist3_dat_o[9] ,
    \wbd_mbist3_dat_o[8] ,
    \wbd_mbist3_dat_o[7] ,
    \wbd_mbist3_dat_o[6] ,
    \wbd_mbist3_dat_o[5] ,
    \wbd_mbist3_dat_o[4] ,
    \wbd_mbist3_dat_o[3] ,
    \wbd_mbist3_dat_o[2] ,
    \wbd_mbist3_dat_o[1] ,
    \wbd_mbist3_dat_o[0] }),
    .s3_wbd_sel_o({\wbd_mbist3_sel_o[3] ,
    \wbd_mbist3_sel_o[2] ,
    \wbd_mbist3_sel_o[1] ,
    \wbd_mbist3_sel_o[0] }),
    .s4_wbd_adr_o({\wbd_mbist4_adr_o[10] ,
    \wbd_mbist4_adr_o[9] ,
    \wbd_mbist4_adr_o[8] ,
    \wbd_mbist4_adr_o[7] ,
    \wbd_mbist4_adr_o[6] ,
    \wbd_mbist4_adr_o[5] ,
    \wbd_mbist4_adr_o[4] ,
    \wbd_mbist4_adr_o[3] ,
    \wbd_mbist4_adr_o[2] ,
    \wbd_mbist4_adr_o[1] ,
    \wbd_mbist4_adr_o[0] }),
    .s4_wbd_dat_i({\wbd_mbist4_dat_i[31] ,
    \wbd_mbist4_dat_i[30] ,
    \wbd_mbist4_dat_i[29] ,
    \wbd_mbist4_dat_i[28] ,
    \wbd_mbist4_dat_i[27] ,
    \wbd_mbist4_dat_i[26] ,
    \wbd_mbist4_dat_i[25] ,
    \wbd_mbist4_dat_i[24] ,
    \wbd_mbist4_dat_i[23] ,
    \wbd_mbist4_dat_i[22] ,
    \wbd_mbist4_dat_i[21] ,
    \wbd_mbist4_dat_i[20] ,
    \wbd_mbist4_dat_i[19] ,
    \wbd_mbist4_dat_i[18] ,
    \wbd_mbist4_dat_i[17] ,
    \wbd_mbist4_dat_i[16] ,
    \wbd_mbist4_dat_i[15] ,
    \wbd_mbist4_dat_i[14] ,
    \wbd_mbist4_dat_i[13] ,
    \wbd_mbist4_dat_i[12] ,
    \wbd_mbist4_dat_i[11] ,
    \wbd_mbist4_dat_i[10] ,
    \wbd_mbist4_dat_i[9] ,
    \wbd_mbist4_dat_i[8] ,
    \wbd_mbist4_dat_i[7] ,
    \wbd_mbist4_dat_i[6] ,
    \wbd_mbist4_dat_i[5] ,
    \wbd_mbist4_dat_i[4] ,
    \wbd_mbist4_dat_i[3] ,
    \wbd_mbist4_dat_i[2] ,
    \wbd_mbist4_dat_i[1] ,
    \wbd_mbist4_dat_i[0] }),
    .s4_wbd_dat_o({\wbd_mbist4_dat_o[31] ,
    \wbd_mbist4_dat_o[30] ,
    \wbd_mbist4_dat_o[29] ,
    \wbd_mbist4_dat_o[28] ,
    \wbd_mbist4_dat_o[27] ,
    \wbd_mbist4_dat_o[26] ,
    \wbd_mbist4_dat_o[25] ,
    \wbd_mbist4_dat_o[24] ,
    \wbd_mbist4_dat_o[23] ,
    \wbd_mbist4_dat_o[22] ,
    \wbd_mbist4_dat_o[21] ,
    \wbd_mbist4_dat_o[20] ,
    \wbd_mbist4_dat_o[19] ,
    \wbd_mbist4_dat_o[18] ,
    \wbd_mbist4_dat_o[17] ,
    \wbd_mbist4_dat_o[16] ,
    \wbd_mbist4_dat_o[15] ,
    \wbd_mbist4_dat_o[14] ,
    \wbd_mbist4_dat_o[13] ,
    \wbd_mbist4_dat_o[12] ,
    \wbd_mbist4_dat_o[11] ,
    \wbd_mbist4_dat_o[10] ,
    \wbd_mbist4_dat_o[9] ,
    \wbd_mbist4_dat_o[8] ,
    \wbd_mbist4_dat_o[7] ,
    \wbd_mbist4_dat_o[6] ,
    \wbd_mbist4_dat_o[5] ,
    \wbd_mbist4_dat_o[4] ,
    \wbd_mbist4_dat_o[3] ,
    \wbd_mbist4_dat_o[2] ,
    \wbd_mbist4_dat_o[1] ,
    \wbd_mbist4_dat_o[0] }),
    .s4_wbd_sel_o({\wbd_mbist4_sel_o[3] ,
    \wbd_mbist4_sel_o[2] ,
    \wbd_mbist4_sel_o[1] ,
    \wbd_mbist4_sel_o[0] }),
    .s5_wbd_adr_o({\wbd_mbist5_adr_o[9] ,
    \wbd_mbist5_adr_o[8] ,
    \wbd_mbist5_adr_o[7] ,
    \wbd_mbist5_adr_o[6] ,
    \wbd_mbist5_adr_o[5] ,
    \wbd_mbist5_adr_o[4] ,
    \wbd_mbist5_adr_o[3] ,
    \wbd_mbist5_adr_o[2] ,
    \wbd_mbist5_adr_o[1] ,
    \wbd_mbist5_adr_o[0] }),
    .s5_wbd_dat_i({\wbd_mbist5_dat_i[31] ,
    \wbd_mbist5_dat_i[30] ,
    \wbd_mbist5_dat_i[29] ,
    \wbd_mbist5_dat_i[28] ,
    \wbd_mbist5_dat_i[27] ,
    \wbd_mbist5_dat_i[26] ,
    \wbd_mbist5_dat_i[25] ,
    \wbd_mbist5_dat_i[24] ,
    \wbd_mbist5_dat_i[23] ,
    \wbd_mbist5_dat_i[22] ,
    \wbd_mbist5_dat_i[21] ,
    \wbd_mbist5_dat_i[20] ,
    \wbd_mbist5_dat_i[19] ,
    \wbd_mbist5_dat_i[18] ,
    \wbd_mbist5_dat_i[17] ,
    \wbd_mbist5_dat_i[16] ,
    \wbd_mbist5_dat_i[15] ,
    \wbd_mbist5_dat_i[14] ,
    \wbd_mbist5_dat_i[13] ,
    \wbd_mbist5_dat_i[12] ,
    \wbd_mbist5_dat_i[11] ,
    \wbd_mbist5_dat_i[10] ,
    \wbd_mbist5_dat_i[9] ,
    \wbd_mbist5_dat_i[8] ,
    \wbd_mbist5_dat_i[7] ,
    \wbd_mbist5_dat_i[6] ,
    \wbd_mbist5_dat_i[5] ,
    \wbd_mbist5_dat_i[4] ,
    \wbd_mbist5_dat_i[3] ,
    \wbd_mbist5_dat_i[2] ,
    \wbd_mbist5_dat_i[1] ,
    \wbd_mbist5_dat_i[0] }),
    .s5_wbd_dat_o({\wbd_mbist5_dat_o[31] ,
    \wbd_mbist5_dat_o[30] ,
    \wbd_mbist5_dat_o[29] ,
    \wbd_mbist5_dat_o[28] ,
    \wbd_mbist5_dat_o[27] ,
    \wbd_mbist5_dat_o[26] ,
    \wbd_mbist5_dat_o[25] ,
    \wbd_mbist5_dat_o[24] ,
    \wbd_mbist5_dat_o[23] ,
    \wbd_mbist5_dat_o[22] ,
    \wbd_mbist5_dat_o[21] ,
    \wbd_mbist5_dat_o[20] ,
    \wbd_mbist5_dat_o[19] ,
    \wbd_mbist5_dat_o[18] ,
    \wbd_mbist5_dat_o[17] ,
    \wbd_mbist5_dat_o[16] ,
    \wbd_mbist5_dat_o[15] ,
    \wbd_mbist5_dat_o[14] ,
    \wbd_mbist5_dat_o[13] ,
    \wbd_mbist5_dat_o[12] ,
    \wbd_mbist5_dat_o[11] ,
    \wbd_mbist5_dat_o[10] ,
    \wbd_mbist5_dat_o[9] ,
    \wbd_mbist5_dat_o[8] ,
    \wbd_mbist5_dat_o[7] ,
    \wbd_mbist5_dat_o[6] ,
    \wbd_mbist5_dat_o[5] ,
    \wbd_mbist5_dat_o[4] ,
    \wbd_mbist5_dat_o[3] ,
    \wbd_mbist5_dat_o[2] ,
    \wbd_mbist5_dat_o[1] ,
    \wbd_mbist5_dat_o[0] }),
    .s5_wbd_sel_o({\wbd_mbist5_sel_o[3] ,
    \wbd_mbist5_sel_o[2] ,
    \wbd_mbist5_sel_o[1] ,
    \wbd_mbist5_sel_o[0] }),
    .s6_wbd_adr_o({\wbd_mbist6_adr_o[9] ,
    \wbd_mbist6_adr_o[8] ,
    \wbd_mbist6_adr_o[7] ,
    \wbd_mbist6_adr_o[6] ,
    \wbd_mbist6_adr_o[5] ,
    \wbd_mbist6_adr_o[4] ,
    \wbd_mbist6_adr_o[3] ,
    \wbd_mbist6_adr_o[2] ,
    \wbd_mbist6_adr_o[1] ,
    \wbd_mbist6_adr_o[0] }),
    .s6_wbd_dat_i({\wbd_mbist6_dat_i[31] ,
    \wbd_mbist6_dat_i[30] ,
    \wbd_mbist6_dat_i[29] ,
    \wbd_mbist6_dat_i[28] ,
    \wbd_mbist6_dat_i[27] ,
    \wbd_mbist6_dat_i[26] ,
    \wbd_mbist6_dat_i[25] ,
    \wbd_mbist6_dat_i[24] ,
    \wbd_mbist6_dat_i[23] ,
    \wbd_mbist6_dat_i[22] ,
    \wbd_mbist6_dat_i[21] ,
    \wbd_mbist6_dat_i[20] ,
    \wbd_mbist6_dat_i[19] ,
    \wbd_mbist6_dat_i[18] ,
    \wbd_mbist6_dat_i[17] ,
    \wbd_mbist6_dat_i[16] ,
    \wbd_mbist6_dat_i[15] ,
    \wbd_mbist6_dat_i[14] ,
    \wbd_mbist6_dat_i[13] ,
    \wbd_mbist6_dat_i[12] ,
    \wbd_mbist6_dat_i[11] ,
    \wbd_mbist6_dat_i[10] ,
    \wbd_mbist6_dat_i[9] ,
    \wbd_mbist6_dat_i[8] ,
    \wbd_mbist6_dat_i[7] ,
    \wbd_mbist6_dat_i[6] ,
    \wbd_mbist6_dat_i[5] ,
    \wbd_mbist6_dat_i[4] ,
    \wbd_mbist6_dat_i[3] ,
    \wbd_mbist6_dat_i[2] ,
    \wbd_mbist6_dat_i[1] ,
    \wbd_mbist6_dat_i[0] }),
    .s6_wbd_dat_o({\wbd_mbist6_dat_o[31] ,
    \wbd_mbist6_dat_o[30] ,
    \wbd_mbist6_dat_o[29] ,
    \wbd_mbist6_dat_o[28] ,
    \wbd_mbist6_dat_o[27] ,
    \wbd_mbist6_dat_o[26] ,
    \wbd_mbist6_dat_o[25] ,
    \wbd_mbist6_dat_o[24] ,
    \wbd_mbist6_dat_o[23] ,
    \wbd_mbist6_dat_o[22] ,
    \wbd_mbist6_dat_o[21] ,
    \wbd_mbist6_dat_o[20] ,
    \wbd_mbist6_dat_o[19] ,
    \wbd_mbist6_dat_o[18] ,
    \wbd_mbist6_dat_o[17] ,
    \wbd_mbist6_dat_o[16] ,
    \wbd_mbist6_dat_o[15] ,
    \wbd_mbist6_dat_o[14] ,
    \wbd_mbist6_dat_o[13] ,
    \wbd_mbist6_dat_o[12] ,
    \wbd_mbist6_dat_o[11] ,
    \wbd_mbist6_dat_o[10] ,
    \wbd_mbist6_dat_o[9] ,
    \wbd_mbist6_dat_o[8] ,
    \wbd_mbist6_dat_o[7] ,
    \wbd_mbist6_dat_o[6] ,
    \wbd_mbist6_dat_o[5] ,
    \wbd_mbist6_dat_o[4] ,
    \wbd_mbist6_dat_o[3] ,
    \wbd_mbist6_dat_o[2] ,
    \wbd_mbist6_dat_o[1] ,
    \wbd_mbist6_dat_o[0] }),
    .s6_wbd_sel_o({\wbd_mbist6_sel_o[3] ,
    \wbd_mbist6_sel_o[2] ,
    \wbd_mbist6_sel_o[1] ,
    \wbd_mbist6_sel_o[0] }),
    .s7_wbd_adr_o({\wbd_mbist7_adr_o[9] ,
    \wbd_mbist7_adr_o[8] ,
    \wbd_mbist7_adr_o[7] ,
    \wbd_mbist7_adr_o[6] ,
    \wbd_mbist7_adr_o[5] ,
    \wbd_mbist7_adr_o[4] ,
    \wbd_mbist7_adr_o[3] ,
    \wbd_mbist7_adr_o[2] ,
    \wbd_mbist7_adr_o[1] ,
    \wbd_mbist7_adr_o[0] }),
    .s7_wbd_dat_i({\wbd_mbist7_dat_i[31] ,
    \wbd_mbist7_dat_i[30] ,
    \wbd_mbist7_dat_i[29] ,
    \wbd_mbist7_dat_i[28] ,
    \wbd_mbist7_dat_i[27] ,
    \wbd_mbist7_dat_i[26] ,
    \wbd_mbist7_dat_i[25] ,
    \wbd_mbist7_dat_i[24] ,
    \wbd_mbist7_dat_i[23] ,
    \wbd_mbist7_dat_i[22] ,
    \wbd_mbist7_dat_i[21] ,
    \wbd_mbist7_dat_i[20] ,
    \wbd_mbist7_dat_i[19] ,
    \wbd_mbist7_dat_i[18] ,
    \wbd_mbist7_dat_i[17] ,
    \wbd_mbist7_dat_i[16] ,
    \wbd_mbist7_dat_i[15] ,
    \wbd_mbist7_dat_i[14] ,
    \wbd_mbist7_dat_i[13] ,
    \wbd_mbist7_dat_i[12] ,
    \wbd_mbist7_dat_i[11] ,
    \wbd_mbist7_dat_i[10] ,
    \wbd_mbist7_dat_i[9] ,
    \wbd_mbist7_dat_i[8] ,
    \wbd_mbist7_dat_i[7] ,
    \wbd_mbist7_dat_i[6] ,
    \wbd_mbist7_dat_i[5] ,
    \wbd_mbist7_dat_i[4] ,
    \wbd_mbist7_dat_i[3] ,
    \wbd_mbist7_dat_i[2] ,
    \wbd_mbist7_dat_i[1] ,
    \wbd_mbist7_dat_i[0] }),
    .s7_wbd_dat_o({\wbd_mbist7_dat_o[31] ,
    \wbd_mbist7_dat_o[30] ,
    \wbd_mbist7_dat_o[29] ,
    \wbd_mbist7_dat_o[28] ,
    \wbd_mbist7_dat_o[27] ,
    \wbd_mbist7_dat_o[26] ,
    \wbd_mbist7_dat_o[25] ,
    \wbd_mbist7_dat_o[24] ,
    \wbd_mbist7_dat_o[23] ,
    \wbd_mbist7_dat_o[22] ,
    \wbd_mbist7_dat_o[21] ,
    \wbd_mbist7_dat_o[20] ,
    \wbd_mbist7_dat_o[19] ,
    \wbd_mbist7_dat_o[18] ,
    \wbd_mbist7_dat_o[17] ,
    \wbd_mbist7_dat_o[16] ,
    \wbd_mbist7_dat_o[15] ,
    \wbd_mbist7_dat_o[14] ,
    \wbd_mbist7_dat_o[13] ,
    \wbd_mbist7_dat_o[12] ,
    \wbd_mbist7_dat_o[11] ,
    \wbd_mbist7_dat_o[10] ,
    \wbd_mbist7_dat_o[9] ,
    \wbd_mbist7_dat_o[8] ,
    \wbd_mbist7_dat_o[7] ,
    \wbd_mbist7_dat_o[6] ,
    \wbd_mbist7_dat_o[5] ,
    \wbd_mbist7_dat_o[4] ,
    \wbd_mbist7_dat_o[3] ,
    \wbd_mbist7_dat_o[2] ,
    \wbd_mbist7_dat_o[1] ,
    \wbd_mbist7_dat_o[0] }),
    .s7_wbd_sel_o({\wbd_mbist7_sel_o[3] ,
    \wbd_mbist7_sel_o[2] ,
    \wbd_mbist7_sel_o[1] ,
    \wbd_mbist7_sel_o[0] }),
    .s8_wbd_adr_o({\wbd_mbist8_adr_o[9] ,
    \wbd_mbist8_adr_o[8] ,
    \wbd_mbist8_adr_o[7] ,
    \wbd_mbist8_adr_o[6] ,
    \wbd_mbist8_adr_o[5] ,
    \wbd_mbist8_adr_o[4] ,
    \wbd_mbist8_adr_o[3] ,
    \wbd_mbist8_adr_o[2] ,
    \wbd_mbist8_adr_o[1] ,
    \wbd_mbist8_adr_o[0] }),
    .s8_wbd_dat_i({\wbd_mbist8_dat_i[31] ,
    \wbd_mbist8_dat_i[30] ,
    \wbd_mbist8_dat_i[29] ,
    \wbd_mbist8_dat_i[28] ,
    \wbd_mbist8_dat_i[27] ,
    \wbd_mbist8_dat_i[26] ,
    \wbd_mbist8_dat_i[25] ,
    \wbd_mbist8_dat_i[24] ,
    \wbd_mbist8_dat_i[23] ,
    \wbd_mbist8_dat_i[22] ,
    \wbd_mbist8_dat_i[21] ,
    \wbd_mbist8_dat_i[20] ,
    \wbd_mbist8_dat_i[19] ,
    \wbd_mbist8_dat_i[18] ,
    \wbd_mbist8_dat_i[17] ,
    \wbd_mbist8_dat_i[16] ,
    \wbd_mbist8_dat_i[15] ,
    \wbd_mbist8_dat_i[14] ,
    \wbd_mbist8_dat_i[13] ,
    \wbd_mbist8_dat_i[12] ,
    \wbd_mbist8_dat_i[11] ,
    \wbd_mbist8_dat_i[10] ,
    \wbd_mbist8_dat_i[9] ,
    \wbd_mbist8_dat_i[8] ,
    \wbd_mbist8_dat_i[7] ,
    \wbd_mbist8_dat_i[6] ,
    \wbd_mbist8_dat_i[5] ,
    \wbd_mbist8_dat_i[4] ,
    \wbd_mbist8_dat_i[3] ,
    \wbd_mbist8_dat_i[2] ,
    \wbd_mbist8_dat_i[1] ,
    \wbd_mbist8_dat_i[0] }),
    .s8_wbd_dat_o({\wbd_mbist8_dat_o[31] ,
    \wbd_mbist8_dat_o[30] ,
    \wbd_mbist8_dat_o[29] ,
    \wbd_mbist8_dat_o[28] ,
    \wbd_mbist8_dat_o[27] ,
    \wbd_mbist8_dat_o[26] ,
    \wbd_mbist8_dat_o[25] ,
    \wbd_mbist8_dat_o[24] ,
    \wbd_mbist8_dat_o[23] ,
    \wbd_mbist8_dat_o[22] ,
    \wbd_mbist8_dat_o[21] ,
    \wbd_mbist8_dat_o[20] ,
    \wbd_mbist8_dat_o[19] ,
    \wbd_mbist8_dat_o[18] ,
    \wbd_mbist8_dat_o[17] ,
    \wbd_mbist8_dat_o[16] ,
    \wbd_mbist8_dat_o[15] ,
    \wbd_mbist8_dat_o[14] ,
    \wbd_mbist8_dat_o[13] ,
    \wbd_mbist8_dat_o[12] ,
    \wbd_mbist8_dat_o[11] ,
    \wbd_mbist8_dat_o[10] ,
    \wbd_mbist8_dat_o[9] ,
    \wbd_mbist8_dat_o[8] ,
    \wbd_mbist8_dat_o[7] ,
    \wbd_mbist8_dat_o[6] ,
    \wbd_mbist8_dat_o[5] ,
    \wbd_mbist8_dat_o[4] ,
    \wbd_mbist8_dat_o[3] ,
    \wbd_mbist8_dat_o[2] ,
    \wbd_mbist8_dat_o[1] ,
    \wbd_mbist8_dat_o[0] }),
    .s8_wbd_sel_o({\wbd_mbist8_sel_o[3] ,
    \wbd_mbist8_sel_o[2] ,
    \wbd_mbist8_sel_o[1] ,
    \wbd_mbist8_sel_o[0] }),
    .scan_si({\scan_out_mbist8[7] ,
    \scan_out_mbist8[6] ,
    \scan_out_mbist8[5] ,
    \scan_out_mbist8[4] ,
    \scan_out_mbist8[3] ,
    \scan_out_mbist8[2] ,
    \scan_out_mbist8[1] ,
    \scan_out_mbist8[0] }),
    .scan_so({\scan_out_wbi[7] ,
    \scan_out_wbi[6] ,
    \scan_out_wbi[5] ,
    \scan_out_wbi[4] ,
    \scan_out_wbi[3] ,
    \scan_out_wbi[2] ,
    \scan_out_wbi[1] ,
    \scan_out_wbi[0] }));
 mbist_top1 u_mbist1 (.bist_correct(\bist_correct[0] ),
    .bist_done(\bist_done[0] ),
    .bist_en(\bist_en_int[0] ),
    .bist_error(\bist_error[0] ),
    .bist_load(\bist_load_int[0] ),
    .bist_run(\bist_run_int[0] ),
    .bist_sdi(\bist_sdi_int[0] ),
    .bist_sdo(\bist_sdo[0] ),
    .bist_shift(\bist_shift_int[0] ),
    .mem_cen_a(mem1_cen_a),
    .mem_cen_b(mem1_cen_b),
    .mem_clk_a(mem1_clk_a),
    .mem_clk_b(mem1_clk_b),
    .mem_web_b(mem1_web_b),
    .rst_n(bist_rst_n),
    .scan_en(scan_en_mbist2),
    .scan_en_o(scan_en_mbist1),
    .scan_mode(scan_mode_mbist2),
    .scan_mode_o(scan_mode_mbist1),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_ack_o(wbd_mbist1_ack_i),
    .wb_clk_i(wbd_clk_mbist1),
    .wb_cyc_i(wbd_mbist1_cyc_o),
    .wb_stb_i(wbd_mbist1_stb_o),
    .wb_we_i(wbd_mbist1_we_o),
    .wbd_clk_int(wbd_clk_mbist1_int),
    .wbd_clk_mbist(wbd_clk_mbist1),
    .bist_error_cnt({\bist_error_cnt0[3] ,
    \bist_error_cnt0[2] ,
    \bist_error_cnt0[1] ,
    \bist_error_cnt0[0] }),
    .cfg_cska_mbist({\cfg_clk_ctrl2[3] ,
    \cfg_clk_ctrl2[2] ,
    \cfg_clk_ctrl2[1] ,
    \cfg_clk_ctrl2[0] }),
    .mem_addr_a({\mem1_addr_a[10] ,
    \mem1_addr_a[9] ,
    \mem1_addr_a[8] ,
    \mem1_addr_a[7] ,
    \mem1_addr_a[6] ,
    \mem1_addr_a[5] ,
    \mem1_addr_a[4] ,
    \mem1_addr_a[3] ,
    \mem1_addr_a[2] }),
    .mem_addr_b({\mem1_addr_b[10] ,
    \mem1_addr_b[9] ,
    \mem1_addr_b[8] ,
    \mem1_addr_b[7] ,
    \mem1_addr_b[6] ,
    \mem1_addr_b[5] ,
    \mem1_addr_b[4] ,
    \mem1_addr_b[3] ,
    \mem1_addr_b[2] }),
    .mem_din_b({\mem1_din_b[31] ,
    \mem1_din_b[30] ,
    \mem1_din_b[29] ,
    \mem1_din_b[28] ,
    \mem1_din_b[27] ,
    \mem1_din_b[26] ,
    \mem1_din_b[25] ,
    \mem1_din_b[24] ,
    \mem1_din_b[23] ,
    \mem1_din_b[22] ,
    \mem1_din_b[21] ,
    \mem1_din_b[20] ,
    \mem1_din_b[19] ,
    \mem1_din_b[18] ,
    \mem1_din_b[17] ,
    \mem1_din_b[16] ,
    \mem1_din_b[15] ,
    \mem1_din_b[14] ,
    \mem1_din_b[13] ,
    \mem1_din_b[12] ,
    \mem1_din_b[11] ,
    \mem1_din_b[10] ,
    \mem1_din_b[9] ,
    \mem1_din_b[8] ,
    \mem1_din_b[7] ,
    \mem1_din_b[6] ,
    \mem1_din_b[5] ,
    \mem1_din_b[4] ,
    \mem1_din_b[3] ,
    \mem1_din_b[2] ,
    \mem1_din_b[1] ,
    \mem1_din_b[0] }),
    .mem_dout_a({\mem1_dout_a[31] ,
    \mem1_dout_a[30] ,
    \mem1_dout_a[29] ,
    \mem1_dout_a[28] ,
    \mem1_dout_a[27] ,
    \mem1_dout_a[26] ,
    \mem1_dout_a[25] ,
    \mem1_dout_a[24] ,
    \mem1_dout_a[23] ,
    \mem1_dout_a[22] ,
    \mem1_dout_a[21] ,
    \mem1_dout_a[20] ,
    \mem1_dout_a[19] ,
    \mem1_dout_a[18] ,
    \mem1_dout_a[17] ,
    \mem1_dout_a[16] ,
    \mem1_dout_a[15] ,
    \mem1_dout_a[14] ,
    \mem1_dout_a[13] ,
    \mem1_dout_a[12] ,
    \mem1_dout_a[11] ,
    \mem1_dout_a[10] ,
    \mem1_dout_a[9] ,
    \mem1_dout_a[8] ,
    \mem1_dout_a[7] ,
    \mem1_dout_a[6] ,
    \mem1_dout_a[5] ,
    \mem1_dout_a[4] ,
    \mem1_dout_a[3] ,
    \mem1_dout_a[2] ,
    \mem1_dout_a[1] ,
    \mem1_dout_a[0] }),
    .mem_mask_b({\mem1_mask_b[3] ,
    \mem1_mask_b[2] ,
    \mem1_mask_b[1] ,
    \mem1_mask_b[0] }),
    .scan_si({\scan_out_mbist2[7] ,
    \scan_out_mbist2[6] ,
    \scan_out_mbist2[5] ,
    \scan_out_mbist2[4] ,
    \scan_out_mbist2[3] ,
    \scan_out_mbist2[2] ,
    \scan_out_mbist2[1] ,
    \scan_out_mbist2[0] }),
    .scan_so({\scan_out_mbist1[7] ,
    \scan_out_mbist1[6] ,
    \scan_out_mbist1[5] ,
    \scan_out_mbist1[4] ,
    \scan_out_mbist1[3] ,
    \scan_out_mbist1[2] ,
    \scan_out_mbist1[1] ,
    \scan_out_mbist1[0] }),
    .wb_adr_i({\wbd_mbist1_adr_o[10] ,
    \wbd_mbist1_adr_o[9] ,
    \wbd_mbist1_adr_o[8] ,
    \wbd_mbist1_adr_o[7] ,
    \wbd_mbist1_adr_o[6] ,
    \wbd_mbist1_adr_o[5] ,
    \wbd_mbist1_adr_o[4] ,
    \wbd_mbist1_adr_o[3] ,
    \wbd_mbist1_adr_o[2] }),
    .wb_dat_i({\wbd_mbist1_dat_o[31] ,
    \wbd_mbist1_dat_o[30] ,
    \wbd_mbist1_dat_o[29] ,
    \wbd_mbist1_dat_o[28] ,
    \wbd_mbist1_dat_o[27] ,
    \wbd_mbist1_dat_o[26] ,
    \wbd_mbist1_dat_o[25] ,
    \wbd_mbist1_dat_o[24] ,
    \wbd_mbist1_dat_o[23] ,
    \wbd_mbist1_dat_o[22] ,
    \wbd_mbist1_dat_o[21] ,
    \wbd_mbist1_dat_o[20] ,
    \wbd_mbist1_dat_o[19] ,
    \wbd_mbist1_dat_o[18] ,
    \wbd_mbist1_dat_o[17] ,
    \wbd_mbist1_dat_o[16] ,
    \wbd_mbist1_dat_o[15] ,
    \wbd_mbist1_dat_o[14] ,
    \wbd_mbist1_dat_o[13] ,
    \wbd_mbist1_dat_o[12] ,
    \wbd_mbist1_dat_o[11] ,
    \wbd_mbist1_dat_o[10] ,
    \wbd_mbist1_dat_o[9] ,
    \wbd_mbist1_dat_o[8] ,
    \wbd_mbist1_dat_o[7] ,
    \wbd_mbist1_dat_o[6] ,
    \wbd_mbist1_dat_o[5] ,
    \wbd_mbist1_dat_o[4] ,
    \wbd_mbist1_dat_o[3] ,
    \wbd_mbist1_dat_o[2] ,
    \wbd_mbist1_dat_o[1] ,
    \wbd_mbist1_dat_o[0] }),
    .wb_dat_o({\wbd_mbist1_dat_i[31] ,
    \wbd_mbist1_dat_i[30] ,
    \wbd_mbist1_dat_i[29] ,
    \wbd_mbist1_dat_i[28] ,
    \wbd_mbist1_dat_i[27] ,
    \wbd_mbist1_dat_i[26] ,
    \wbd_mbist1_dat_i[25] ,
    \wbd_mbist1_dat_i[24] ,
    \wbd_mbist1_dat_i[23] ,
    \wbd_mbist1_dat_i[22] ,
    \wbd_mbist1_dat_i[21] ,
    \wbd_mbist1_dat_i[20] ,
    \wbd_mbist1_dat_i[19] ,
    \wbd_mbist1_dat_i[18] ,
    \wbd_mbist1_dat_i[17] ,
    \wbd_mbist1_dat_i[16] ,
    \wbd_mbist1_dat_i[15] ,
    \wbd_mbist1_dat_i[14] ,
    \wbd_mbist1_dat_i[13] ,
    \wbd_mbist1_dat_i[12] ,
    \wbd_mbist1_dat_i[11] ,
    \wbd_mbist1_dat_i[10] ,
    \wbd_mbist1_dat_i[9] ,
    \wbd_mbist1_dat_i[8] ,
    \wbd_mbist1_dat_i[7] ,
    \wbd_mbist1_dat_i[6] ,
    \wbd_mbist1_dat_i[5] ,
    \wbd_mbist1_dat_i[4] ,
    \wbd_mbist1_dat_i[3] ,
    \wbd_mbist1_dat_i[2] ,
    \wbd_mbist1_dat_i[1] ,
    \wbd_mbist1_dat_i[0] }),
    .wb_sel_i({\wbd_mbist1_sel_o[3] ,
    \wbd_mbist1_sel_o[2] ,
    \wbd_mbist1_sel_o[1] ,
    \wbd_mbist1_sel_o[0] }));
 mbist_top1 u_mbist2 (.bist_correct(\bist_correct[1] ),
    .bist_done(\bist_done[1] ),
    .bist_en(\bist_en_int[1] ),
    .bist_error(\bist_error[1] ),
    .bist_load(\bist_load_int[1] ),
    .bist_run(\bist_run_int[1] ),
    .bist_sdi(\bist_sdi_int[1] ),
    .bist_sdo(\bist_sdo[1] ),
    .bist_shift(\bist_shift_int[1] ),
    .mem_cen_a(mem2_cen_a),
    .mem_cen_b(mem2_cen_b),
    .mem_clk_a(mem2_clk_a),
    .mem_clk_b(mem2_clk_b),
    .mem_web_b(mem2_web_b),
    .rst_n(bist_rst_n),
    .scan_en(scan_en_mbist3),
    .scan_en_o(scan_en_mbist2),
    .scan_mode(scan_mode_mbist3),
    .scan_mode_o(scan_mode_mbist2),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_ack_o(wbd_mbist2_ack_i),
    .wb_clk_i(wbd_clk_mbist2),
    .wb_cyc_i(wbd_mbist2_cyc_o),
    .wb_stb_i(wbd_mbist2_stb_o),
    .wb_we_i(wbd_mbist2_we_o),
    .wbd_clk_int(wbd_clk_mbist2_int),
    .wbd_clk_mbist(wbd_clk_mbist2),
    .bist_error_cnt({\bist_error_cnt1[3] ,
    \bist_error_cnt1[2] ,
    \bist_error_cnt1[1] ,
    \bist_error_cnt1[0] }),
    .cfg_cska_mbist({\cfg_clk_ctrl2[7] ,
    \cfg_clk_ctrl2[6] ,
    \cfg_clk_ctrl2[5] ,
    \cfg_clk_ctrl2[4] }),
    .mem_addr_a({\mem2_addr_a[10] ,
    \mem2_addr_a[9] ,
    \mem2_addr_a[8] ,
    \mem2_addr_a[7] ,
    \mem2_addr_a[6] ,
    \mem2_addr_a[5] ,
    \mem2_addr_a[4] ,
    \mem2_addr_a[3] ,
    \mem2_addr_a[2] }),
    .mem_addr_b({\mem2_addr_b[10] ,
    \mem2_addr_b[9] ,
    \mem2_addr_b[8] ,
    \mem2_addr_b[7] ,
    \mem2_addr_b[6] ,
    \mem2_addr_b[5] ,
    \mem2_addr_b[4] ,
    \mem2_addr_b[3] ,
    \mem2_addr_b[2] }),
    .mem_din_b({\mem2_din_b[31] ,
    \mem2_din_b[30] ,
    \mem2_din_b[29] ,
    \mem2_din_b[28] ,
    \mem2_din_b[27] ,
    \mem2_din_b[26] ,
    \mem2_din_b[25] ,
    \mem2_din_b[24] ,
    \mem2_din_b[23] ,
    \mem2_din_b[22] ,
    \mem2_din_b[21] ,
    \mem2_din_b[20] ,
    \mem2_din_b[19] ,
    \mem2_din_b[18] ,
    \mem2_din_b[17] ,
    \mem2_din_b[16] ,
    \mem2_din_b[15] ,
    \mem2_din_b[14] ,
    \mem2_din_b[13] ,
    \mem2_din_b[12] ,
    \mem2_din_b[11] ,
    \mem2_din_b[10] ,
    \mem2_din_b[9] ,
    \mem2_din_b[8] ,
    \mem2_din_b[7] ,
    \mem2_din_b[6] ,
    \mem2_din_b[5] ,
    \mem2_din_b[4] ,
    \mem2_din_b[3] ,
    \mem2_din_b[2] ,
    \mem2_din_b[1] ,
    \mem2_din_b[0] }),
    .mem_dout_a({\mem2_dout_a[31] ,
    \mem2_dout_a[30] ,
    \mem2_dout_a[29] ,
    \mem2_dout_a[28] ,
    \mem2_dout_a[27] ,
    \mem2_dout_a[26] ,
    \mem2_dout_a[25] ,
    \mem2_dout_a[24] ,
    \mem2_dout_a[23] ,
    \mem2_dout_a[22] ,
    \mem2_dout_a[21] ,
    \mem2_dout_a[20] ,
    \mem2_dout_a[19] ,
    \mem2_dout_a[18] ,
    \mem2_dout_a[17] ,
    \mem2_dout_a[16] ,
    \mem2_dout_a[15] ,
    \mem2_dout_a[14] ,
    \mem2_dout_a[13] ,
    \mem2_dout_a[12] ,
    \mem2_dout_a[11] ,
    \mem2_dout_a[10] ,
    \mem2_dout_a[9] ,
    \mem2_dout_a[8] ,
    \mem2_dout_a[7] ,
    \mem2_dout_a[6] ,
    \mem2_dout_a[5] ,
    \mem2_dout_a[4] ,
    \mem2_dout_a[3] ,
    \mem2_dout_a[2] ,
    \mem2_dout_a[1] ,
    \mem2_dout_a[0] }),
    .mem_mask_b({\mem2_mask_b[3] ,
    \mem2_mask_b[2] ,
    \mem2_mask_b[1] ,
    \mem2_mask_b[0] }),
    .scan_si({\scan_out_mbist3[7] ,
    \scan_out_mbist3[6] ,
    \scan_out_mbist3[5] ,
    \scan_out_mbist3[4] ,
    \scan_out_mbist3[3] ,
    \scan_out_mbist3[2] ,
    \scan_out_mbist3[1] ,
    \scan_out_mbist3[0] }),
    .scan_so({\scan_out_mbist2[7] ,
    \scan_out_mbist2[6] ,
    \scan_out_mbist2[5] ,
    \scan_out_mbist2[4] ,
    \scan_out_mbist2[3] ,
    \scan_out_mbist2[2] ,
    \scan_out_mbist2[1] ,
    \scan_out_mbist2[0] }),
    .wb_adr_i({\wbd_mbist2_adr_o[10] ,
    \wbd_mbist2_adr_o[9] ,
    \wbd_mbist2_adr_o[8] ,
    \wbd_mbist2_adr_o[7] ,
    \wbd_mbist2_adr_o[6] ,
    \wbd_mbist2_adr_o[5] ,
    \wbd_mbist2_adr_o[4] ,
    \wbd_mbist2_adr_o[3] ,
    \wbd_mbist2_adr_o[2] }),
    .wb_dat_i({\wbd_mbist2_dat_o[31] ,
    \wbd_mbist2_dat_o[30] ,
    \wbd_mbist2_dat_o[29] ,
    \wbd_mbist2_dat_o[28] ,
    \wbd_mbist2_dat_o[27] ,
    \wbd_mbist2_dat_o[26] ,
    \wbd_mbist2_dat_o[25] ,
    \wbd_mbist2_dat_o[24] ,
    \wbd_mbist2_dat_o[23] ,
    \wbd_mbist2_dat_o[22] ,
    \wbd_mbist2_dat_o[21] ,
    \wbd_mbist2_dat_o[20] ,
    \wbd_mbist2_dat_o[19] ,
    \wbd_mbist2_dat_o[18] ,
    \wbd_mbist2_dat_o[17] ,
    \wbd_mbist2_dat_o[16] ,
    \wbd_mbist2_dat_o[15] ,
    \wbd_mbist2_dat_o[14] ,
    \wbd_mbist2_dat_o[13] ,
    \wbd_mbist2_dat_o[12] ,
    \wbd_mbist2_dat_o[11] ,
    \wbd_mbist2_dat_o[10] ,
    \wbd_mbist2_dat_o[9] ,
    \wbd_mbist2_dat_o[8] ,
    \wbd_mbist2_dat_o[7] ,
    \wbd_mbist2_dat_o[6] ,
    \wbd_mbist2_dat_o[5] ,
    \wbd_mbist2_dat_o[4] ,
    \wbd_mbist2_dat_o[3] ,
    \wbd_mbist2_dat_o[2] ,
    \wbd_mbist2_dat_o[1] ,
    \wbd_mbist2_dat_o[0] }),
    .wb_dat_o({\wbd_mbist2_dat_i[31] ,
    \wbd_mbist2_dat_i[30] ,
    \wbd_mbist2_dat_i[29] ,
    \wbd_mbist2_dat_i[28] ,
    \wbd_mbist2_dat_i[27] ,
    \wbd_mbist2_dat_i[26] ,
    \wbd_mbist2_dat_i[25] ,
    \wbd_mbist2_dat_i[24] ,
    \wbd_mbist2_dat_i[23] ,
    \wbd_mbist2_dat_i[22] ,
    \wbd_mbist2_dat_i[21] ,
    \wbd_mbist2_dat_i[20] ,
    \wbd_mbist2_dat_i[19] ,
    \wbd_mbist2_dat_i[18] ,
    \wbd_mbist2_dat_i[17] ,
    \wbd_mbist2_dat_i[16] ,
    \wbd_mbist2_dat_i[15] ,
    \wbd_mbist2_dat_i[14] ,
    \wbd_mbist2_dat_i[13] ,
    \wbd_mbist2_dat_i[12] ,
    \wbd_mbist2_dat_i[11] ,
    \wbd_mbist2_dat_i[10] ,
    \wbd_mbist2_dat_i[9] ,
    \wbd_mbist2_dat_i[8] ,
    \wbd_mbist2_dat_i[7] ,
    \wbd_mbist2_dat_i[6] ,
    \wbd_mbist2_dat_i[5] ,
    \wbd_mbist2_dat_i[4] ,
    \wbd_mbist2_dat_i[3] ,
    \wbd_mbist2_dat_i[2] ,
    \wbd_mbist2_dat_i[1] ,
    \wbd_mbist2_dat_i[0] }),
    .wb_sel_i({\wbd_mbist2_sel_o[3] ,
    \wbd_mbist2_sel_o[2] ,
    \wbd_mbist2_sel_o[1] ,
    \wbd_mbist2_sel_o[0] }));
 mbist_top1 u_mbist3 (.bist_correct(\bist_correct[2] ),
    .bist_done(\bist_done[2] ),
    .bist_en(\bist_en_int[2] ),
    .bist_error(\bist_error[2] ),
    .bist_load(\bist_load_int[2] ),
    .bist_run(\bist_run_int[2] ),
    .bist_sdi(\bist_sdi_int[2] ),
    .bist_sdo(\bist_sdo[2] ),
    .bist_shift(\bist_shift_int[2] ),
    .mem_cen_a(mem3_cen_a),
    .mem_cen_b(mem3_cen_b),
    .mem_clk_a(mem3_clk_a),
    .mem_clk_b(mem3_clk_b),
    .mem_web_b(mem3_web_b),
    .rst_n(bist_rst_n),
    .scan_en(scan_en_mbist4),
    .scan_en_o(scan_en_mbist3),
    .scan_mode(scan_mode_mbist4),
    .scan_mode_o(scan_mode_mbist3),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_ack_o(wbd_mbist3_ack_i),
    .wb_clk_i(wbd_clk_mbist3),
    .wb_cyc_i(wbd_mbist3_cyc_o),
    .wb_stb_i(wbd_mbist3_stb_o),
    .wb_we_i(wbd_mbist3_we_o),
    .wbd_clk_int(wbd_clk_mbist3_int),
    .wbd_clk_mbist(wbd_clk_mbist3),
    .bist_error_cnt({\bist_error_cnt2[3] ,
    \bist_error_cnt2[2] ,
    \bist_error_cnt2[1] ,
    \bist_error_cnt2[0] }),
    .cfg_cska_mbist({\cfg_clk_ctrl2[11] ,
    \cfg_clk_ctrl2[10] ,
    \cfg_clk_ctrl2[9] ,
    \cfg_clk_ctrl2[8] }),
    .mem_addr_a({\mem3_addr_a[10] ,
    \mem3_addr_a[9] ,
    \mem3_addr_a[8] ,
    \mem3_addr_a[7] ,
    \mem3_addr_a[6] ,
    \mem3_addr_a[5] ,
    \mem3_addr_a[4] ,
    \mem3_addr_a[3] ,
    \mem3_addr_a[2] }),
    .mem_addr_b({\mem3_addr_b[10] ,
    \mem3_addr_b[9] ,
    \mem3_addr_b[8] ,
    \mem3_addr_b[7] ,
    \mem3_addr_b[6] ,
    \mem3_addr_b[5] ,
    \mem3_addr_b[4] ,
    \mem3_addr_b[3] ,
    \mem3_addr_b[2] }),
    .mem_din_b({\mem3_din_b[31] ,
    \mem3_din_b[30] ,
    \mem3_din_b[29] ,
    \mem3_din_b[28] ,
    \mem3_din_b[27] ,
    \mem3_din_b[26] ,
    \mem3_din_b[25] ,
    \mem3_din_b[24] ,
    \mem3_din_b[23] ,
    \mem3_din_b[22] ,
    \mem3_din_b[21] ,
    \mem3_din_b[20] ,
    \mem3_din_b[19] ,
    \mem3_din_b[18] ,
    \mem3_din_b[17] ,
    \mem3_din_b[16] ,
    \mem3_din_b[15] ,
    \mem3_din_b[14] ,
    \mem3_din_b[13] ,
    \mem3_din_b[12] ,
    \mem3_din_b[11] ,
    \mem3_din_b[10] ,
    \mem3_din_b[9] ,
    \mem3_din_b[8] ,
    \mem3_din_b[7] ,
    \mem3_din_b[6] ,
    \mem3_din_b[5] ,
    \mem3_din_b[4] ,
    \mem3_din_b[3] ,
    \mem3_din_b[2] ,
    \mem3_din_b[1] ,
    \mem3_din_b[0] }),
    .mem_dout_a({\mem3_dout_a[31] ,
    \mem3_dout_a[30] ,
    \mem3_dout_a[29] ,
    \mem3_dout_a[28] ,
    \mem3_dout_a[27] ,
    \mem3_dout_a[26] ,
    \mem3_dout_a[25] ,
    \mem3_dout_a[24] ,
    \mem3_dout_a[23] ,
    \mem3_dout_a[22] ,
    \mem3_dout_a[21] ,
    \mem3_dout_a[20] ,
    \mem3_dout_a[19] ,
    \mem3_dout_a[18] ,
    \mem3_dout_a[17] ,
    \mem3_dout_a[16] ,
    \mem3_dout_a[15] ,
    \mem3_dout_a[14] ,
    \mem3_dout_a[13] ,
    \mem3_dout_a[12] ,
    \mem3_dout_a[11] ,
    \mem3_dout_a[10] ,
    \mem3_dout_a[9] ,
    \mem3_dout_a[8] ,
    \mem3_dout_a[7] ,
    \mem3_dout_a[6] ,
    \mem3_dout_a[5] ,
    \mem3_dout_a[4] ,
    \mem3_dout_a[3] ,
    \mem3_dout_a[2] ,
    \mem3_dout_a[1] ,
    \mem3_dout_a[0] }),
    .mem_mask_b({\mem3_mask_b[3] ,
    \mem3_mask_b[2] ,
    \mem3_mask_b[1] ,
    \mem3_mask_b[0] }),
    .scan_si({\scan_out_mbist4[7] ,
    \scan_out_mbist4[6] ,
    \scan_out_mbist4[5] ,
    \scan_out_mbist4[4] ,
    \scan_out_mbist4[3] ,
    \scan_out_mbist4[2] ,
    \scan_out_mbist4[1] ,
    \scan_out_mbist4[0] }),
    .scan_so({\scan_out_mbist3[7] ,
    \scan_out_mbist3[6] ,
    \scan_out_mbist3[5] ,
    \scan_out_mbist3[4] ,
    \scan_out_mbist3[3] ,
    \scan_out_mbist3[2] ,
    \scan_out_mbist3[1] ,
    \scan_out_mbist3[0] }),
    .wb_adr_i({\wbd_mbist3_adr_o[10] ,
    \wbd_mbist3_adr_o[9] ,
    \wbd_mbist3_adr_o[8] ,
    \wbd_mbist3_adr_o[7] ,
    \wbd_mbist3_adr_o[6] ,
    \wbd_mbist3_adr_o[5] ,
    \wbd_mbist3_adr_o[4] ,
    \wbd_mbist3_adr_o[3] ,
    \wbd_mbist3_adr_o[2] }),
    .wb_dat_i({\wbd_mbist3_dat_o[31] ,
    \wbd_mbist3_dat_o[30] ,
    \wbd_mbist3_dat_o[29] ,
    \wbd_mbist3_dat_o[28] ,
    \wbd_mbist3_dat_o[27] ,
    \wbd_mbist3_dat_o[26] ,
    \wbd_mbist3_dat_o[25] ,
    \wbd_mbist3_dat_o[24] ,
    \wbd_mbist3_dat_o[23] ,
    \wbd_mbist3_dat_o[22] ,
    \wbd_mbist3_dat_o[21] ,
    \wbd_mbist3_dat_o[20] ,
    \wbd_mbist3_dat_o[19] ,
    \wbd_mbist3_dat_o[18] ,
    \wbd_mbist3_dat_o[17] ,
    \wbd_mbist3_dat_o[16] ,
    \wbd_mbist3_dat_o[15] ,
    \wbd_mbist3_dat_o[14] ,
    \wbd_mbist3_dat_o[13] ,
    \wbd_mbist3_dat_o[12] ,
    \wbd_mbist3_dat_o[11] ,
    \wbd_mbist3_dat_o[10] ,
    \wbd_mbist3_dat_o[9] ,
    \wbd_mbist3_dat_o[8] ,
    \wbd_mbist3_dat_o[7] ,
    \wbd_mbist3_dat_o[6] ,
    \wbd_mbist3_dat_o[5] ,
    \wbd_mbist3_dat_o[4] ,
    \wbd_mbist3_dat_o[3] ,
    \wbd_mbist3_dat_o[2] ,
    \wbd_mbist3_dat_o[1] ,
    \wbd_mbist3_dat_o[0] }),
    .wb_dat_o({\wbd_mbist3_dat_i[31] ,
    \wbd_mbist3_dat_i[30] ,
    \wbd_mbist3_dat_i[29] ,
    \wbd_mbist3_dat_i[28] ,
    \wbd_mbist3_dat_i[27] ,
    \wbd_mbist3_dat_i[26] ,
    \wbd_mbist3_dat_i[25] ,
    \wbd_mbist3_dat_i[24] ,
    \wbd_mbist3_dat_i[23] ,
    \wbd_mbist3_dat_i[22] ,
    \wbd_mbist3_dat_i[21] ,
    \wbd_mbist3_dat_i[20] ,
    \wbd_mbist3_dat_i[19] ,
    \wbd_mbist3_dat_i[18] ,
    \wbd_mbist3_dat_i[17] ,
    \wbd_mbist3_dat_i[16] ,
    \wbd_mbist3_dat_i[15] ,
    \wbd_mbist3_dat_i[14] ,
    \wbd_mbist3_dat_i[13] ,
    \wbd_mbist3_dat_i[12] ,
    \wbd_mbist3_dat_i[11] ,
    \wbd_mbist3_dat_i[10] ,
    \wbd_mbist3_dat_i[9] ,
    \wbd_mbist3_dat_i[8] ,
    \wbd_mbist3_dat_i[7] ,
    \wbd_mbist3_dat_i[6] ,
    \wbd_mbist3_dat_i[5] ,
    \wbd_mbist3_dat_i[4] ,
    \wbd_mbist3_dat_i[3] ,
    \wbd_mbist3_dat_i[2] ,
    \wbd_mbist3_dat_i[1] ,
    \wbd_mbist3_dat_i[0] }),
    .wb_sel_i({\wbd_mbist3_sel_o[3] ,
    \wbd_mbist3_sel_o[2] ,
    \wbd_mbist3_sel_o[1] ,
    \wbd_mbist3_sel_o[0] }));
 mbist_top1 u_mbist4 (.bist_correct(\bist_correct[3] ),
    .bist_done(\bist_done[3] ),
    .bist_en(\bist_en_int[3] ),
    .bist_error(\bist_error[3] ),
    .bist_load(\bist_load_int[3] ),
    .bist_run(\bist_run_int[3] ),
    .bist_sdi(\bist_sdi_int[3] ),
    .bist_sdo(\bist_sdo[3] ),
    .bist_shift(\bist_shift_int[3] ),
    .mem_cen_a(mem4_cen_a),
    .mem_cen_b(mem4_cen_b),
    .mem_clk_a(mem4_clk_a),
    .mem_clk_b(mem4_clk_b),
    .mem_web_b(mem4_web_b),
    .rst_n(bist_rst_n),
    .scan_en(scan_en_wbi),
    .scan_en_o(scan_en_mbist4),
    .scan_mode(scan_mode_wbi),
    .scan_mode_o(scan_mode_mbist4),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_ack_o(wbd_mbist4_ack_i),
    .wb_clk_i(wbd_clk_mbist4),
    .wb_cyc_i(wbd_mbist4_cyc_o),
    .wb_stb_i(wbd_mbist4_stb_o),
    .wb_we_i(wbd_mbist4_we_o),
    .wbd_clk_int(wbd_clk_mbist4_int),
    .wbd_clk_mbist(wbd_clk_mbist4),
    .bist_error_cnt({\bist_error_cnt3[3] ,
    \bist_error_cnt3[2] ,
    \bist_error_cnt3[1] ,
    \bist_error_cnt3[0] }),
    .cfg_cska_mbist({\cfg_clk_ctrl2[15] ,
    \cfg_clk_ctrl2[14] ,
    \cfg_clk_ctrl2[13] ,
    \cfg_clk_ctrl2[12] }),
    .mem_addr_a({\mem4_addr_a[10] ,
    \mem4_addr_a[9] ,
    \mem4_addr_a[8] ,
    \mem4_addr_a[7] ,
    \mem4_addr_a[6] ,
    \mem4_addr_a[5] ,
    \mem4_addr_a[4] ,
    \mem4_addr_a[3] ,
    \mem4_addr_a[2] }),
    .mem_addr_b({\mem4_addr_b[10] ,
    \mem4_addr_b[9] ,
    \mem4_addr_b[8] ,
    \mem4_addr_b[7] ,
    \mem4_addr_b[6] ,
    \mem4_addr_b[5] ,
    \mem4_addr_b[4] ,
    \mem4_addr_b[3] ,
    \mem4_addr_b[2] }),
    .mem_din_b({\mem4_din_b[31] ,
    \mem4_din_b[30] ,
    \mem4_din_b[29] ,
    \mem4_din_b[28] ,
    \mem4_din_b[27] ,
    \mem4_din_b[26] ,
    \mem4_din_b[25] ,
    \mem4_din_b[24] ,
    \mem4_din_b[23] ,
    \mem4_din_b[22] ,
    \mem4_din_b[21] ,
    \mem4_din_b[20] ,
    \mem4_din_b[19] ,
    \mem4_din_b[18] ,
    \mem4_din_b[17] ,
    \mem4_din_b[16] ,
    \mem4_din_b[15] ,
    \mem4_din_b[14] ,
    \mem4_din_b[13] ,
    \mem4_din_b[12] ,
    \mem4_din_b[11] ,
    \mem4_din_b[10] ,
    \mem4_din_b[9] ,
    \mem4_din_b[8] ,
    \mem4_din_b[7] ,
    \mem4_din_b[6] ,
    \mem4_din_b[5] ,
    \mem4_din_b[4] ,
    \mem4_din_b[3] ,
    \mem4_din_b[2] ,
    \mem4_din_b[1] ,
    \mem4_din_b[0] }),
    .mem_dout_a({\mem4_dout_a[31] ,
    \mem4_dout_a[30] ,
    \mem4_dout_a[29] ,
    \mem4_dout_a[28] ,
    \mem4_dout_a[27] ,
    \mem4_dout_a[26] ,
    \mem4_dout_a[25] ,
    \mem4_dout_a[24] ,
    \mem4_dout_a[23] ,
    \mem4_dout_a[22] ,
    \mem4_dout_a[21] ,
    \mem4_dout_a[20] ,
    \mem4_dout_a[19] ,
    \mem4_dout_a[18] ,
    \mem4_dout_a[17] ,
    \mem4_dout_a[16] ,
    \mem4_dout_a[15] ,
    \mem4_dout_a[14] ,
    \mem4_dout_a[13] ,
    \mem4_dout_a[12] ,
    \mem4_dout_a[11] ,
    \mem4_dout_a[10] ,
    \mem4_dout_a[9] ,
    \mem4_dout_a[8] ,
    \mem4_dout_a[7] ,
    \mem4_dout_a[6] ,
    \mem4_dout_a[5] ,
    \mem4_dout_a[4] ,
    \mem4_dout_a[3] ,
    \mem4_dout_a[2] ,
    \mem4_dout_a[1] ,
    \mem4_dout_a[0] }),
    .mem_mask_b({\mem4_mask_b[3] ,
    \mem4_mask_b[2] ,
    \mem4_mask_b[1] ,
    \mem4_mask_b[0] }),
    .scan_si({\scan_out_wbi[7] ,
    \scan_out_wbi[6] ,
    \scan_out_wbi[5] ,
    \scan_out_wbi[4] ,
    \scan_out_wbi[3] ,
    \scan_out_wbi[2] ,
    \scan_out_wbi[1] ,
    \scan_out_wbi[0] }),
    .scan_so({\scan_out_mbist4[7] ,
    \scan_out_mbist4[6] ,
    \scan_out_mbist4[5] ,
    \scan_out_mbist4[4] ,
    \scan_out_mbist4[3] ,
    \scan_out_mbist4[2] ,
    \scan_out_mbist4[1] ,
    \scan_out_mbist4[0] }),
    .wb_adr_i({\wbd_mbist4_adr_o[10] ,
    \wbd_mbist4_adr_o[9] ,
    \wbd_mbist4_adr_o[8] ,
    \wbd_mbist4_adr_o[7] ,
    \wbd_mbist4_adr_o[6] ,
    \wbd_mbist4_adr_o[5] ,
    \wbd_mbist4_adr_o[4] ,
    \wbd_mbist4_adr_o[3] ,
    \wbd_mbist4_adr_o[2] }),
    .wb_dat_i({\wbd_mbist4_dat_o[31] ,
    \wbd_mbist4_dat_o[30] ,
    \wbd_mbist4_dat_o[29] ,
    \wbd_mbist4_dat_o[28] ,
    \wbd_mbist4_dat_o[27] ,
    \wbd_mbist4_dat_o[26] ,
    \wbd_mbist4_dat_o[25] ,
    \wbd_mbist4_dat_o[24] ,
    \wbd_mbist4_dat_o[23] ,
    \wbd_mbist4_dat_o[22] ,
    \wbd_mbist4_dat_o[21] ,
    \wbd_mbist4_dat_o[20] ,
    \wbd_mbist4_dat_o[19] ,
    \wbd_mbist4_dat_o[18] ,
    \wbd_mbist4_dat_o[17] ,
    \wbd_mbist4_dat_o[16] ,
    \wbd_mbist4_dat_o[15] ,
    \wbd_mbist4_dat_o[14] ,
    \wbd_mbist4_dat_o[13] ,
    \wbd_mbist4_dat_o[12] ,
    \wbd_mbist4_dat_o[11] ,
    \wbd_mbist4_dat_o[10] ,
    \wbd_mbist4_dat_o[9] ,
    \wbd_mbist4_dat_o[8] ,
    \wbd_mbist4_dat_o[7] ,
    \wbd_mbist4_dat_o[6] ,
    \wbd_mbist4_dat_o[5] ,
    \wbd_mbist4_dat_o[4] ,
    \wbd_mbist4_dat_o[3] ,
    \wbd_mbist4_dat_o[2] ,
    \wbd_mbist4_dat_o[1] ,
    \wbd_mbist4_dat_o[0] }),
    .wb_dat_o({\wbd_mbist4_dat_i[31] ,
    \wbd_mbist4_dat_i[30] ,
    \wbd_mbist4_dat_i[29] ,
    \wbd_mbist4_dat_i[28] ,
    \wbd_mbist4_dat_i[27] ,
    \wbd_mbist4_dat_i[26] ,
    \wbd_mbist4_dat_i[25] ,
    \wbd_mbist4_dat_i[24] ,
    \wbd_mbist4_dat_i[23] ,
    \wbd_mbist4_dat_i[22] ,
    \wbd_mbist4_dat_i[21] ,
    \wbd_mbist4_dat_i[20] ,
    \wbd_mbist4_dat_i[19] ,
    \wbd_mbist4_dat_i[18] ,
    \wbd_mbist4_dat_i[17] ,
    \wbd_mbist4_dat_i[16] ,
    \wbd_mbist4_dat_i[15] ,
    \wbd_mbist4_dat_i[14] ,
    \wbd_mbist4_dat_i[13] ,
    \wbd_mbist4_dat_i[12] ,
    \wbd_mbist4_dat_i[11] ,
    \wbd_mbist4_dat_i[10] ,
    \wbd_mbist4_dat_i[9] ,
    \wbd_mbist4_dat_i[8] ,
    \wbd_mbist4_dat_i[7] ,
    \wbd_mbist4_dat_i[6] ,
    \wbd_mbist4_dat_i[5] ,
    \wbd_mbist4_dat_i[4] ,
    \wbd_mbist4_dat_i[3] ,
    \wbd_mbist4_dat_i[2] ,
    \wbd_mbist4_dat_i[1] ,
    \wbd_mbist4_dat_i[0] }),
    .wb_sel_i({\wbd_mbist4_sel_o[3] ,
    \wbd_mbist4_sel_o[2] ,
    \wbd_mbist4_sel_o[1] ,
    \wbd_mbist4_sel_o[0] }));
 mbist_top2 u_mbist5 (.bist_correct(\bist_correct[4] ),
    .bist_done(\bist_done[4] ),
    .bist_en(\bist_en_int[4] ),
    .bist_error(\bist_error[4] ),
    .bist_load(\bist_load_int[4] ),
    .bist_run(\bist_run_int[4] ),
    .bist_sdi(\bist_sdi_int[4] ),
    .bist_sdo(\bist_sdo[4] ),
    .bist_shift(\bist_shift_int[4] ),
    .mem_cen_a(mem5_cen_a),
    .mem_cen_b(mem5_cen_b),
    .mem_clk_a(mem5_clk_a),
    .mem_clk_b(mem5_clk_b),
    .mem_web_b(mem5_web_b),
    .rst_n(bist_rst_n),
    .scan_en(scan_en_glbl),
    .scan_en_o(scan_en_mbist5),
    .scan_mode(scan_mode_glbl),
    .scan_mode_o(scan_mode_mbist5),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_ack_o(wbd_mbist5_ack_i),
    .wb_clk_i(wbd_clk_mbist5),
    .wb_cyc_i(wbd_mbist5_cyc_o),
    .wb_stb_i(wbd_mbist5_stb_o),
    .wb_we_i(wbd_mbist5_we_o),
    .wbd_clk_int(wbd_clk_mbist5_int),
    .wbd_clk_mbist(wbd_clk_mbist5),
    .bist_error_cnt({\bist_error_cnt4[3] ,
    \bist_error_cnt4[2] ,
    \bist_error_cnt4[1] ,
    \bist_error_cnt4[0] }),
    .cfg_cska_mbist({\cfg_clk_ctrl2[19] ,
    \cfg_clk_ctrl2[18] ,
    \cfg_clk_ctrl2[17] ,
    \cfg_clk_ctrl2[16] }),
    .mem_addr_a({\mem5_addr_a[9] ,
    \mem5_addr_a[8] ,
    \mem5_addr_a[7] ,
    \mem5_addr_a[6] ,
    \mem5_addr_a[5] ,
    \mem5_addr_a[4] ,
    \mem5_addr_a[3] ,
    \mem5_addr_a[2] }),
    .mem_addr_b({\mem5_addr_b[9] ,
    \mem5_addr_b[8] ,
    \mem5_addr_b[7] ,
    \mem5_addr_b[6] ,
    \mem5_addr_b[5] ,
    \mem5_addr_b[4] ,
    \mem5_addr_b[3] ,
    \mem5_addr_b[2] }),
    .mem_din_b({\mem5_din_b[31] ,
    \mem5_din_b[30] ,
    \mem5_din_b[29] ,
    \mem5_din_b[28] ,
    \mem5_din_b[27] ,
    \mem5_din_b[26] ,
    \mem5_din_b[25] ,
    \mem5_din_b[24] ,
    \mem5_din_b[23] ,
    \mem5_din_b[22] ,
    \mem5_din_b[21] ,
    \mem5_din_b[20] ,
    \mem5_din_b[19] ,
    \mem5_din_b[18] ,
    \mem5_din_b[17] ,
    \mem5_din_b[16] ,
    \mem5_din_b[15] ,
    \mem5_din_b[14] ,
    \mem5_din_b[13] ,
    \mem5_din_b[12] ,
    \mem5_din_b[11] ,
    \mem5_din_b[10] ,
    \mem5_din_b[9] ,
    \mem5_din_b[8] ,
    \mem5_din_b[7] ,
    \mem5_din_b[6] ,
    \mem5_din_b[5] ,
    \mem5_din_b[4] ,
    \mem5_din_b[3] ,
    \mem5_din_b[2] ,
    \mem5_din_b[1] ,
    \mem5_din_b[0] }),
    .mem_dout_a({\mem5_dout_a[31] ,
    \mem5_dout_a[30] ,
    \mem5_dout_a[29] ,
    \mem5_dout_a[28] ,
    \mem5_dout_a[27] ,
    \mem5_dout_a[26] ,
    \mem5_dout_a[25] ,
    \mem5_dout_a[24] ,
    \mem5_dout_a[23] ,
    \mem5_dout_a[22] ,
    \mem5_dout_a[21] ,
    \mem5_dout_a[20] ,
    \mem5_dout_a[19] ,
    \mem5_dout_a[18] ,
    \mem5_dout_a[17] ,
    \mem5_dout_a[16] ,
    \mem5_dout_a[15] ,
    \mem5_dout_a[14] ,
    \mem5_dout_a[13] ,
    \mem5_dout_a[12] ,
    \mem5_dout_a[11] ,
    \mem5_dout_a[10] ,
    \mem5_dout_a[9] ,
    \mem5_dout_a[8] ,
    \mem5_dout_a[7] ,
    \mem5_dout_a[6] ,
    \mem5_dout_a[5] ,
    \mem5_dout_a[4] ,
    \mem5_dout_a[3] ,
    \mem5_dout_a[2] ,
    \mem5_dout_a[1] ,
    \mem5_dout_a[0] }),
    .mem_mask_b({\mem5_mask_b[3] ,
    \mem5_mask_b[2] ,
    \mem5_mask_b[1] ,
    \mem5_mask_b[0] }),
    .scan_si({\scan_out_glbl[7] ,
    \scan_out_glbl[6] ,
    \scan_out_glbl[5] ,
    \scan_out_glbl[4] ,
    \scan_out_glbl[3] ,
    \scan_out_glbl[2] ,
    \scan_out_glbl[1] ,
    \scan_out_glbl[0] }),
    .scan_so({\scan_out_mbist5[7] ,
    \scan_out_mbist5[6] ,
    \scan_out_mbist5[5] ,
    \scan_out_mbist5[4] ,
    \scan_out_mbist5[3] ,
    \scan_out_mbist5[2] ,
    \scan_out_mbist5[1] ,
    \scan_out_mbist5[0] }),
    .wb_adr_i({\wbd_mbist5_adr_o[9] ,
    \wbd_mbist5_adr_o[8] ,
    \wbd_mbist5_adr_o[7] ,
    \wbd_mbist5_adr_o[6] ,
    \wbd_mbist5_adr_o[5] ,
    \wbd_mbist5_adr_o[4] ,
    \wbd_mbist5_adr_o[3] ,
    \wbd_mbist5_adr_o[2] }),
    .wb_dat_i({\wbd_mbist5_dat_o[31] ,
    \wbd_mbist5_dat_o[30] ,
    \wbd_mbist5_dat_o[29] ,
    \wbd_mbist5_dat_o[28] ,
    \wbd_mbist5_dat_o[27] ,
    \wbd_mbist5_dat_o[26] ,
    \wbd_mbist5_dat_o[25] ,
    \wbd_mbist5_dat_o[24] ,
    \wbd_mbist5_dat_o[23] ,
    \wbd_mbist5_dat_o[22] ,
    \wbd_mbist5_dat_o[21] ,
    \wbd_mbist5_dat_o[20] ,
    \wbd_mbist5_dat_o[19] ,
    \wbd_mbist5_dat_o[18] ,
    \wbd_mbist5_dat_o[17] ,
    \wbd_mbist5_dat_o[16] ,
    \wbd_mbist5_dat_o[15] ,
    \wbd_mbist5_dat_o[14] ,
    \wbd_mbist5_dat_o[13] ,
    \wbd_mbist5_dat_o[12] ,
    \wbd_mbist5_dat_o[11] ,
    \wbd_mbist5_dat_o[10] ,
    \wbd_mbist5_dat_o[9] ,
    \wbd_mbist5_dat_o[8] ,
    \wbd_mbist5_dat_o[7] ,
    \wbd_mbist5_dat_o[6] ,
    \wbd_mbist5_dat_o[5] ,
    \wbd_mbist5_dat_o[4] ,
    \wbd_mbist5_dat_o[3] ,
    \wbd_mbist5_dat_o[2] ,
    \wbd_mbist5_dat_o[1] ,
    \wbd_mbist5_dat_o[0] }),
    .wb_dat_o({\wbd_mbist5_dat_i[31] ,
    \wbd_mbist5_dat_i[30] ,
    \wbd_mbist5_dat_i[29] ,
    \wbd_mbist5_dat_i[28] ,
    \wbd_mbist5_dat_i[27] ,
    \wbd_mbist5_dat_i[26] ,
    \wbd_mbist5_dat_i[25] ,
    \wbd_mbist5_dat_i[24] ,
    \wbd_mbist5_dat_i[23] ,
    \wbd_mbist5_dat_i[22] ,
    \wbd_mbist5_dat_i[21] ,
    \wbd_mbist5_dat_i[20] ,
    \wbd_mbist5_dat_i[19] ,
    \wbd_mbist5_dat_i[18] ,
    \wbd_mbist5_dat_i[17] ,
    \wbd_mbist5_dat_i[16] ,
    \wbd_mbist5_dat_i[15] ,
    \wbd_mbist5_dat_i[14] ,
    \wbd_mbist5_dat_i[13] ,
    \wbd_mbist5_dat_i[12] ,
    \wbd_mbist5_dat_i[11] ,
    \wbd_mbist5_dat_i[10] ,
    \wbd_mbist5_dat_i[9] ,
    \wbd_mbist5_dat_i[8] ,
    \wbd_mbist5_dat_i[7] ,
    \wbd_mbist5_dat_i[6] ,
    \wbd_mbist5_dat_i[5] ,
    \wbd_mbist5_dat_i[4] ,
    \wbd_mbist5_dat_i[3] ,
    \wbd_mbist5_dat_i[2] ,
    \wbd_mbist5_dat_i[1] ,
    \wbd_mbist5_dat_i[0] }),
    .wb_sel_i({\wbd_mbist5_sel_o[3] ,
    \wbd_mbist5_sel_o[2] ,
    \wbd_mbist5_sel_o[1] ,
    \wbd_mbist5_sel_o[0] }));
 mbist_top2 u_mbist6 (.bist_correct(\bist_correct[5] ),
    .bist_done(\bist_done[5] ),
    .bist_en(\bist_en_int[5] ),
    .bist_error(\bist_error[5] ),
    .bist_load(\bist_load_int[5] ),
    .bist_run(\bist_run_int[5] ),
    .bist_sdi(\bist_sdi_int[5] ),
    .bist_sdo(\bist_sdo[5] ),
    .bist_shift(\bist_shift_int[5] ),
    .mem_cen_a(mem6_cen_a),
    .mem_cen_b(mem6_cen_b),
    .mem_clk_a(mem6_clk_a),
    .mem_clk_b(mem6_clk_b),
    .mem_web_b(mem6_web_b),
    .rst_n(bist_rst_n),
    .scan_en(scan_en_mbist5),
    .scan_en_o(scan_en_mbist6),
    .scan_mode(scan_mode_mbist5),
    .scan_mode_o(scan_mode_mbist6),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_ack_o(wbd_mbist6_ack_i),
    .wb_clk_i(wbd_clk_mbist6),
    .wb_cyc_i(wbd_mbist6_cyc_o),
    .wb_stb_i(wbd_mbist6_stb_o),
    .wb_we_i(wbd_mbist6_we_o),
    .wbd_clk_int(wbd_clk_mbist6_int),
    .wbd_clk_mbist(wbd_clk_mbist6),
    .bist_error_cnt({\bist_error_cnt5[3] ,
    \bist_error_cnt5[2] ,
    \bist_error_cnt5[1] ,
    \bist_error_cnt5[0] }),
    .cfg_cska_mbist({\cfg_clk_ctrl2[23] ,
    \cfg_clk_ctrl2[22] ,
    \cfg_clk_ctrl2[21] ,
    \cfg_clk_ctrl2[20] }),
    .mem_addr_a({\mem6_addr_a[9] ,
    \mem6_addr_a[8] ,
    \mem6_addr_a[7] ,
    \mem6_addr_a[6] ,
    \mem6_addr_a[5] ,
    \mem6_addr_a[4] ,
    \mem6_addr_a[3] ,
    \mem6_addr_a[2] }),
    .mem_addr_b({\mem6_addr_b[9] ,
    \mem6_addr_b[8] ,
    \mem6_addr_b[7] ,
    \mem6_addr_b[6] ,
    \mem6_addr_b[5] ,
    \mem6_addr_b[4] ,
    \mem6_addr_b[3] ,
    \mem6_addr_b[2] }),
    .mem_din_b({\mem6_din_b[31] ,
    \mem6_din_b[30] ,
    \mem6_din_b[29] ,
    \mem6_din_b[28] ,
    \mem6_din_b[27] ,
    \mem6_din_b[26] ,
    \mem6_din_b[25] ,
    \mem6_din_b[24] ,
    \mem6_din_b[23] ,
    \mem6_din_b[22] ,
    \mem6_din_b[21] ,
    \mem6_din_b[20] ,
    \mem6_din_b[19] ,
    \mem6_din_b[18] ,
    \mem6_din_b[17] ,
    \mem6_din_b[16] ,
    \mem6_din_b[15] ,
    \mem6_din_b[14] ,
    \mem6_din_b[13] ,
    \mem6_din_b[12] ,
    \mem6_din_b[11] ,
    \mem6_din_b[10] ,
    \mem6_din_b[9] ,
    \mem6_din_b[8] ,
    \mem6_din_b[7] ,
    \mem6_din_b[6] ,
    \mem6_din_b[5] ,
    \mem6_din_b[4] ,
    \mem6_din_b[3] ,
    \mem6_din_b[2] ,
    \mem6_din_b[1] ,
    \mem6_din_b[0] }),
    .mem_dout_a({\mem6_dout_a[31] ,
    \mem6_dout_a[30] ,
    \mem6_dout_a[29] ,
    \mem6_dout_a[28] ,
    \mem6_dout_a[27] ,
    \mem6_dout_a[26] ,
    \mem6_dout_a[25] ,
    \mem6_dout_a[24] ,
    \mem6_dout_a[23] ,
    \mem6_dout_a[22] ,
    \mem6_dout_a[21] ,
    \mem6_dout_a[20] ,
    \mem6_dout_a[19] ,
    \mem6_dout_a[18] ,
    \mem6_dout_a[17] ,
    \mem6_dout_a[16] ,
    \mem6_dout_a[15] ,
    \mem6_dout_a[14] ,
    \mem6_dout_a[13] ,
    \mem6_dout_a[12] ,
    \mem6_dout_a[11] ,
    \mem6_dout_a[10] ,
    \mem6_dout_a[9] ,
    \mem6_dout_a[8] ,
    \mem6_dout_a[7] ,
    \mem6_dout_a[6] ,
    \mem6_dout_a[5] ,
    \mem6_dout_a[4] ,
    \mem6_dout_a[3] ,
    \mem6_dout_a[2] ,
    \mem6_dout_a[1] ,
    \mem6_dout_a[0] }),
    .mem_mask_b({\mem6_mask_b[3] ,
    \mem6_mask_b[2] ,
    \mem6_mask_b[1] ,
    \mem6_mask_b[0] }),
    .scan_si({\scan_out_mbist5[7] ,
    \scan_out_mbist5[6] ,
    \scan_out_mbist5[5] ,
    \scan_out_mbist5[4] ,
    \scan_out_mbist5[3] ,
    \scan_out_mbist5[2] ,
    \scan_out_mbist5[1] ,
    \scan_out_mbist5[0] }),
    .scan_so({\scan_out_mbist6[7] ,
    \scan_out_mbist6[6] ,
    \scan_out_mbist6[5] ,
    \scan_out_mbist6[4] ,
    \scan_out_mbist6[3] ,
    \scan_out_mbist6[2] ,
    \scan_out_mbist6[1] ,
    \scan_out_mbist6[0] }),
    .wb_adr_i({\wbd_mbist6_adr_o[9] ,
    \wbd_mbist6_adr_o[8] ,
    \wbd_mbist6_adr_o[7] ,
    \wbd_mbist6_adr_o[6] ,
    \wbd_mbist6_adr_o[5] ,
    \wbd_mbist6_adr_o[4] ,
    \wbd_mbist6_adr_o[3] ,
    \wbd_mbist6_adr_o[2] }),
    .wb_dat_i({\wbd_mbist6_dat_o[31] ,
    \wbd_mbist6_dat_o[30] ,
    \wbd_mbist6_dat_o[29] ,
    \wbd_mbist6_dat_o[28] ,
    \wbd_mbist6_dat_o[27] ,
    \wbd_mbist6_dat_o[26] ,
    \wbd_mbist6_dat_o[25] ,
    \wbd_mbist6_dat_o[24] ,
    \wbd_mbist6_dat_o[23] ,
    \wbd_mbist6_dat_o[22] ,
    \wbd_mbist6_dat_o[21] ,
    \wbd_mbist6_dat_o[20] ,
    \wbd_mbist6_dat_o[19] ,
    \wbd_mbist6_dat_o[18] ,
    \wbd_mbist6_dat_o[17] ,
    \wbd_mbist6_dat_o[16] ,
    \wbd_mbist6_dat_o[15] ,
    \wbd_mbist6_dat_o[14] ,
    \wbd_mbist6_dat_o[13] ,
    \wbd_mbist6_dat_o[12] ,
    \wbd_mbist6_dat_o[11] ,
    \wbd_mbist6_dat_o[10] ,
    \wbd_mbist6_dat_o[9] ,
    \wbd_mbist6_dat_o[8] ,
    \wbd_mbist6_dat_o[7] ,
    \wbd_mbist6_dat_o[6] ,
    \wbd_mbist6_dat_o[5] ,
    \wbd_mbist6_dat_o[4] ,
    \wbd_mbist6_dat_o[3] ,
    \wbd_mbist6_dat_o[2] ,
    \wbd_mbist6_dat_o[1] ,
    \wbd_mbist6_dat_o[0] }),
    .wb_dat_o({\wbd_mbist6_dat_i[31] ,
    \wbd_mbist6_dat_i[30] ,
    \wbd_mbist6_dat_i[29] ,
    \wbd_mbist6_dat_i[28] ,
    \wbd_mbist6_dat_i[27] ,
    \wbd_mbist6_dat_i[26] ,
    \wbd_mbist6_dat_i[25] ,
    \wbd_mbist6_dat_i[24] ,
    \wbd_mbist6_dat_i[23] ,
    \wbd_mbist6_dat_i[22] ,
    \wbd_mbist6_dat_i[21] ,
    \wbd_mbist6_dat_i[20] ,
    \wbd_mbist6_dat_i[19] ,
    \wbd_mbist6_dat_i[18] ,
    \wbd_mbist6_dat_i[17] ,
    \wbd_mbist6_dat_i[16] ,
    \wbd_mbist6_dat_i[15] ,
    \wbd_mbist6_dat_i[14] ,
    \wbd_mbist6_dat_i[13] ,
    \wbd_mbist6_dat_i[12] ,
    \wbd_mbist6_dat_i[11] ,
    \wbd_mbist6_dat_i[10] ,
    \wbd_mbist6_dat_i[9] ,
    \wbd_mbist6_dat_i[8] ,
    \wbd_mbist6_dat_i[7] ,
    \wbd_mbist6_dat_i[6] ,
    \wbd_mbist6_dat_i[5] ,
    \wbd_mbist6_dat_i[4] ,
    \wbd_mbist6_dat_i[3] ,
    \wbd_mbist6_dat_i[2] ,
    \wbd_mbist6_dat_i[1] ,
    \wbd_mbist6_dat_i[0] }),
    .wb_sel_i({\wbd_mbist6_sel_o[3] ,
    \wbd_mbist6_sel_o[2] ,
    \wbd_mbist6_sel_o[1] ,
    \wbd_mbist6_sel_o[0] }));
 mbist_top2 u_mbist7 (.bist_correct(\bist_correct[6] ),
    .bist_done(\bist_done[6] ),
    .bist_en(\bist_en_int[6] ),
    .bist_error(\bist_error[6] ),
    .bist_load(\bist_load_int[6] ),
    .bist_run(\bist_run_int[6] ),
    .bist_sdi(\bist_sdi_int[6] ),
    .bist_sdo(\bist_sdo[6] ),
    .bist_shift(\bist_shift_int[6] ),
    .mem_cen_a(mem7_cen_a),
    .mem_cen_b(mem7_cen_b),
    .mem_clk_a(mem7_clk_a),
    .mem_clk_b(mem7_clk_b),
    .mem_web_b(mem7_web_b),
    .rst_n(bist_rst_n),
    .scan_en(scan_en_mbist6),
    .scan_en_o(scan_en_mbist7),
    .scan_mode(scan_mode_mbist6),
    .scan_mode_o(scan_mode_mbist7),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_ack_o(wbd_mbist7_ack_i),
    .wb_clk_i(wbd_clk_mbist7),
    .wb_cyc_i(wbd_mbist7_cyc_o),
    .wb_stb_i(wbd_mbist7_stb_o),
    .wb_we_i(wbd_mbist7_we_o),
    .wbd_clk_int(wbd_clk_mbist7_int),
    .wbd_clk_mbist(wbd_clk_mbist7),
    .bist_error_cnt({\bist_error_cnt6[3] ,
    \bist_error_cnt6[2] ,
    \bist_error_cnt6[1] ,
    \bist_error_cnt6[0] }),
    .cfg_cska_mbist({\cfg_clk_ctrl2[27] ,
    \cfg_clk_ctrl2[26] ,
    \cfg_clk_ctrl2[25] ,
    \cfg_clk_ctrl2[24] }),
    .mem_addr_a({\mem7_addr_a[9] ,
    \mem7_addr_a[8] ,
    \mem7_addr_a[7] ,
    \mem7_addr_a[6] ,
    \mem7_addr_a[5] ,
    \mem7_addr_a[4] ,
    \mem7_addr_a[3] ,
    \mem7_addr_a[2] }),
    .mem_addr_b({\mem7_addr_b[9] ,
    \mem7_addr_b[8] ,
    \mem7_addr_b[7] ,
    \mem7_addr_b[6] ,
    \mem7_addr_b[5] ,
    \mem7_addr_b[4] ,
    \mem7_addr_b[3] ,
    \mem7_addr_b[2] }),
    .mem_din_b({\mem7_din_b[31] ,
    \mem7_din_b[30] ,
    \mem7_din_b[29] ,
    \mem7_din_b[28] ,
    \mem7_din_b[27] ,
    \mem7_din_b[26] ,
    \mem7_din_b[25] ,
    \mem7_din_b[24] ,
    \mem7_din_b[23] ,
    \mem7_din_b[22] ,
    \mem7_din_b[21] ,
    \mem7_din_b[20] ,
    \mem7_din_b[19] ,
    \mem7_din_b[18] ,
    \mem7_din_b[17] ,
    \mem7_din_b[16] ,
    \mem7_din_b[15] ,
    \mem7_din_b[14] ,
    \mem7_din_b[13] ,
    \mem7_din_b[12] ,
    \mem7_din_b[11] ,
    \mem7_din_b[10] ,
    \mem7_din_b[9] ,
    \mem7_din_b[8] ,
    \mem7_din_b[7] ,
    \mem7_din_b[6] ,
    \mem7_din_b[5] ,
    \mem7_din_b[4] ,
    \mem7_din_b[3] ,
    \mem7_din_b[2] ,
    \mem7_din_b[1] ,
    \mem7_din_b[0] }),
    .mem_dout_a({\mem7_dout_a[31] ,
    \mem7_dout_a[30] ,
    \mem7_dout_a[29] ,
    \mem7_dout_a[28] ,
    \mem7_dout_a[27] ,
    \mem7_dout_a[26] ,
    \mem7_dout_a[25] ,
    \mem7_dout_a[24] ,
    \mem7_dout_a[23] ,
    \mem7_dout_a[22] ,
    \mem7_dout_a[21] ,
    \mem7_dout_a[20] ,
    \mem7_dout_a[19] ,
    \mem7_dout_a[18] ,
    \mem7_dout_a[17] ,
    \mem7_dout_a[16] ,
    \mem7_dout_a[15] ,
    \mem7_dout_a[14] ,
    \mem7_dout_a[13] ,
    \mem7_dout_a[12] ,
    \mem7_dout_a[11] ,
    \mem7_dout_a[10] ,
    \mem7_dout_a[9] ,
    \mem7_dout_a[8] ,
    \mem7_dout_a[7] ,
    \mem7_dout_a[6] ,
    \mem7_dout_a[5] ,
    \mem7_dout_a[4] ,
    \mem7_dout_a[3] ,
    \mem7_dout_a[2] ,
    \mem7_dout_a[1] ,
    \mem7_dout_a[0] }),
    .mem_mask_b({\mem7_mask_b[3] ,
    \mem7_mask_b[2] ,
    \mem7_mask_b[1] ,
    \mem7_mask_b[0] }),
    .scan_si({\scan_out_mbist6[7] ,
    \scan_out_mbist6[6] ,
    \scan_out_mbist6[5] ,
    \scan_out_mbist6[4] ,
    \scan_out_mbist6[3] ,
    \scan_out_mbist6[2] ,
    \scan_out_mbist6[1] ,
    \scan_out_mbist6[0] }),
    .scan_so({\scan_out_mbist7[7] ,
    \scan_out_mbist7[6] ,
    \scan_out_mbist7[5] ,
    \scan_out_mbist7[4] ,
    \scan_out_mbist7[3] ,
    \scan_out_mbist7[2] ,
    \scan_out_mbist7[1] ,
    \scan_out_mbist7[0] }),
    .wb_adr_i({\wbd_mbist7_adr_o[9] ,
    \wbd_mbist7_adr_o[8] ,
    \wbd_mbist7_adr_o[7] ,
    \wbd_mbist7_adr_o[6] ,
    \wbd_mbist7_adr_o[5] ,
    \wbd_mbist7_adr_o[4] ,
    \wbd_mbist7_adr_o[3] ,
    \wbd_mbist7_adr_o[2] }),
    .wb_dat_i({\wbd_mbist7_dat_o[31] ,
    \wbd_mbist7_dat_o[30] ,
    \wbd_mbist7_dat_o[29] ,
    \wbd_mbist7_dat_o[28] ,
    \wbd_mbist7_dat_o[27] ,
    \wbd_mbist7_dat_o[26] ,
    \wbd_mbist7_dat_o[25] ,
    \wbd_mbist7_dat_o[24] ,
    \wbd_mbist7_dat_o[23] ,
    \wbd_mbist7_dat_o[22] ,
    \wbd_mbist7_dat_o[21] ,
    \wbd_mbist7_dat_o[20] ,
    \wbd_mbist7_dat_o[19] ,
    \wbd_mbist7_dat_o[18] ,
    \wbd_mbist7_dat_o[17] ,
    \wbd_mbist7_dat_o[16] ,
    \wbd_mbist7_dat_o[15] ,
    \wbd_mbist7_dat_o[14] ,
    \wbd_mbist7_dat_o[13] ,
    \wbd_mbist7_dat_o[12] ,
    \wbd_mbist7_dat_o[11] ,
    \wbd_mbist7_dat_o[10] ,
    \wbd_mbist7_dat_o[9] ,
    \wbd_mbist7_dat_o[8] ,
    \wbd_mbist7_dat_o[7] ,
    \wbd_mbist7_dat_o[6] ,
    \wbd_mbist7_dat_o[5] ,
    \wbd_mbist7_dat_o[4] ,
    \wbd_mbist7_dat_o[3] ,
    \wbd_mbist7_dat_o[2] ,
    \wbd_mbist7_dat_o[1] ,
    \wbd_mbist7_dat_o[0] }),
    .wb_dat_o({\wbd_mbist7_dat_i[31] ,
    \wbd_mbist7_dat_i[30] ,
    \wbd_mbist7_dat_i[29] ,
    \wbd_mbist7_dat_i[28] ,
    \wbd_mbist7_dat_i[27] ,
    \wbd_mbist7_dat_i[26] ,
    \wbd_mbist7_dat_i[25] ,
    \wbd_mbist7_dat_i[24] ,
    \wbd_mbist7_dat_i[23] ,
    \wbd_mbist7_dat_i[22] ,
    \wbd_mbist7_dat_i[21] ,
    \wbd_mbist7_dat_i[20] ,
    \wbd_mbist7_dat_i[19] ,
    \wbd_mbist7_dat_i[18] ,
    \wbd_mbist7_dat_i[17] ,
    \wbd_mbist7_dat_i[16] ,
    \wbd_mbist7_dat_i[15] ,
    \wbd_mbist7_dat_i[14] ,
    \wbd_mbist7_dat_i[13] ,
    \wbd_mbist7_dat_i[12] ,
    \wbd_mbist7_dat_i[11] ,
    \wbd_mbist7_dat_i[10] ,
    \wbd_mbist7_dat_i[9] ,
    \wbd_mbist7_dat_i[8] ,
    \wbd_mbist7_dat_i[7] ,
    \wbd_mbist7_dat_i[6] ,
    \wbd_mbist7_dat_i[5] ,
    \wbd_mbist7_dat_i[4] ,
    \wbd_mbist7_dat_i[3] ,
    \wbd_mbist7_dat_i[2] ,
    \wbd_mbist7_dat_i[1] ,
    \wbd_mbist7_dat_i[0] }),
    .wb_sel_i({\wbd_mbist7_sel_o[3] ,
    \wbd_mbist7_sel_o[2] ,
    \wbd_mbist7_sel_o[1] ,
    \wbd_mbist7_sel_o[0] }));
 mbist_top2 u_mbist8 (.bist_correct(\bist_correct[7] ),
    .bist_done(\bist_done[7] ),
    .bist_en(\bist_en_int[7] ),
    .bist_error(\bist_error[7] ),
    .bist_load(\bist_load_int[7] ),
    .bist_run(\bist_run_int[7] ),
    .bist_sdi(\bist_sdi_int[7] ),
    .bist_sdo(\bist_sdo[7] ),
    .bist_shift(\bist_shift_int[7] ),
    .mem_cen_a(mem8_cen_a),
    .mem_cen_b(mem8_cen_b),
    .mem_clk_a(mem8_clk_a),
    .mem_clk_b(mem8_clk_b),
    .mem_web_b(mem8_web_b),
    .rst_n(bist_rst_n),
    .scan_en(scan_en_mbist7),
    .scan_en_o(scan_en_mbist8),
    .scan_mode(scan_mode_mbist7),
    .scan_mode_o(scan_mode_mbist8),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_ack_o(wbd_mbist8_ack_i),
    .wb_clk_i(wbd_clk_mbist8),
    .wb_cyc_i(wbd_mbist8_cyc_o),
    .wb_stb_i(wbd_mbist8_stb_o),
    .wb_we_i(wbd_mbist8_we_o),
    .wbd_clk_int(wbd_clk_mbist8_int),
    .wbd_clk_mbist(wbd_clk_mbist8),
    .bist_error_cnt({\bist_error_cnt7[3] ,
    \bist_error_cnt7[2] ,
    \bist_error_cnt7[1] ,
    \bist_error_cnt7[0] }),
    .cfg_cska_mbist({\cfg_clk_ctrl2[31] ,
    \cfg_clk_ctrl2[30] ,
    \cfg_clk_ctrl2[29] ,
    \cfg_clk_ctrl2[28] }),
    .mem_addr_a({\mem8_addr_a[9] ,
    \mem8_addr_a[8] ,
    \mem8_addr_a[7] ,
    \mem8_addr_a[6] ,
    \mem8_addr_a[5] ,
    \mem8_addr_a[4] ,
    \mem8_addr_a[3] ,
    \mem8_addr_a[2] }),
    .mem_addr_b({\mem8_addr_b[9] ,
    \mem8_addr_b[8] ,
    \mem8_addr_b[7] ,
    \mem8_addr_b[6] ,
    \mem8_addr_b[5] ,
    \mem8_addr_b[4] ,
    \mem8_addr_b[3] ,
    \mem8_addr_b[2] }),
    .mem_din_b({\mem8_din_b[31] ,
    \mem8_din_b[30] ,
    \mem8_din_b[29] ,
    \mem8_din_b[28] ,
    \mem8_din_b[27] ,
    \mem8_din_b[26] ,
    \mem8_din_b[25] ,
    \mem8_din_b[24] ,
    \mem8_din_b[23] ,
    \mem8_din_b[22] ,
    \mem8_din_b[21] ,
    \mem8_din_b[20] ,
    \mem8_din_b[19] ,
    \mem8_din_b[18] ,
    \mem8_din_b[17] ,
    \mem8_din_b[16] ,
    \mem8_din_b[15] ,
    \mem8_din_b[14] ,
    \mem8_din_b[13] ,
    \mem8_din_b[12] ,
    \mem8_din_b[11] ,
    \mem8_din_b[10] ,
    \mem8_din_b[9] ,
    \mem8_din_b[8] ,
    \mem8_din_b[7] ,
    \mem8_din_b[6] ,
    \mem8_din_b[5] ,
    \mem8_din_b[4] ,
    \mem8_din_b[3] ,
    \mem8_din_b[2] ,
    \mem8_din_b[1] ,
    \mem8_din_b[0] }),
    .mem_dout_a({\mem8_dout_a[31] ,
    \mem8_dout_a[30] ,
    \mem8_dout_a[29] ,
    \mem8_dout_a[28] ,
    \mem8_dout_a[27] ,
    \mem8_dout_a[26] ,
    \mem8_dout_a[25] ,
    \mem8_dout_a[24] ,
    \mem8_dout_a[23] ,
    \mem8_dout_a[22] ,
    \mem8_dout_a[21] ,
    \mem8_dout_a[20] ,
    \mem8_dout_a[19] ,
    \mem8_dout_a[18] ,
    \mem8_dout_a[17] ,
    \mem8_dout_a[16] ,
    \mem8_dout_a[15] ,
    \mem8_dout_a[14] ,
    \mem8_dout_a[13] ,
    \mem8_dout_a[12] ,
    \mem8_dout_a[11] ,
    \mem8_dout_a[10] ,
    \mem8_dout_a[9] ,
    \mem8_dout_a[8] ,
    \mem8_dout_a[7] ,
    \mem8_dout_a[6] ,
    \mem8_dout_a[5] ,
    \mem8_dout_a[4] ,
    \mem8_dout_a[3] ,
    \mem8_dout_a[2] ,
    \mem8_dout_a[1] ,
    \mem8_dout_a[0] }),
    .mem_mask_b({\mem8_mask_b[3] ,
    \mem8_mask_b[2] ,
    \mem8_mask_b[1] ,
    \mem8_mask_b[0] }),
    .scan_si({\scan_out_mbist7[7] ,
    \scan_out_mbist7[6] ,
    \scan_out_mbist7[5] ,
    \scan_out_mbist7[4] ,
    \scan_out_mbist7[3] ,
    \scan_out_mbist7[2] ,
    \scan_out_mbist7[1] ,
    \scan_out_mbist7[0] }),
    .scan_so({\scan_out_mbist8[7] ,
    \scan_out_mbist8[6] ,
    \scan_out_mbist8[5] ,
    \scan_out_mbist8[4] ,
    \scan_out_mbist8[3] ,
    \scan_out_mbist8[2] ,
    \scan_out_mbist8[1] ,
    \scan_out_mbist8[0] }),
    .wb_adr_i({\wbd_mbist8_adr_o[9] ,
    \wbd_mbist8_adr_o[8] ,
    \wbd_mbist8_adr_o[7] ,
    \wbd_mbist8_adr_o[6] ,
    \wbd_mbist8_adr_o[5] ,
    \wbd_mbist8_adr_o[4] ,
    \wbd_mbist8_adr_o[3] ,
    \wbd_mbist8_adr_o[2] }),
    .wb_dat_i({\wbd_mbist8_dat_o[31] ,
    \wbd_mbist8_dat_o[30] ,
    \wbd_mbist8_dat_o[29] ,
    \wbd_mbist8_dat_o[28] ,
    \wbd_mbist8_dat_o[27] ,
    \wbd_mbist8_dat_o[26] ,
    \wbd_mbist8_dat_o[25] ,
    \wbd_mbist8_dat_o[24] ,
    \wbd_mbist8_dat_o[23] ,
    \wbd_mbist8_dat_o[22] ,
    \wbd_mbist8_dat_o[21] ,
    \wbd_mbist8_dat_o[20] ,
    \wbd_mbist8_dat_o[19] ,
    \wbd_mbist8_dat_o[18] ,
    \wbd_mbist8_dat_o[17] ,
    \wbd_mbist8_dat_o[16] ,
    \wbd_mbist8_dat_o[15] ,
    \wbd_mbist8_dat_o[14] ,
    \wbd_mbist8_dat_o[13] ,
    \wbd_mbist8_dat_o[12] ,
    \wbd_mbist8_dat_o[11] ,
    \wbd_mbist8_dat_o[10] ,
    \wbd_mbist8_dat_o[9] ,
    \wbd_mbist8_dat_o[8] ,
    \wbd_mbist8_dat_o[7] ,
    \wbd_mbist8_dat_o[6] ,
    \wbd_mbist8_dat_o[5] ,
    \wbd_mbist8_dat_o[4] ,
    \wbd_mbist8_dat_o[3] ,
    \wbd_mbist8_dat_o[2] ,
    \wbd_mbist8_dat_o[1] ,
    \wbd_mbist8_dat_o[0] }),
    .wb_dat_o({\wbd_mbist8_dat_i[31] ,
    \wbd_mbist8_dat_i[30] ,
    \wbd_mbist8_dat_i[29] ,
    \wbd_mbist8_dat_i[28] ,
    \wbd_mbist8_dat_i[27] ,
    \wbd_mbist8_dat_i[26] ,
    \wbd_mbist8_dat_i[25] ,
    \wbd_mbist8_dat_i[24] ,
    \wbd_mbist8_dat_i[23] ,
    \wbd_mbist8_dat_i[22] ,
    \wbd_mbist8_dat_i[21] ,
    \wbd_mbist8_dat_i[20] ,
    \wbd_mbist8_dat_i[19] ,
    \wbd_mbist8_dat_i[18] ,
    \wbd_mbist8_dat_i[17] ,
    \wbd_mbist8_dat_i[16] ,
    \wbd_mbist8_dat_i[15] ,
    \wbd_mbist8_dat_i[14] ,
    \wbd_mbist8_dat_i[13] ,
    \wbd_mbist8_dat_i[12] ,
    \wbd_mbist8_dat_i[11] ,
    \wbd_mbist8_dat_i[10] ,
    \wbd_mbist8_dat_i[9] ,
    \wbd_mbist8_dat_i[8] ,
    \wbd_mbist8_dat_i[7] ,
    \wbd_mbist8_dat_i[6] ,
    \wbd_mbist8_dat_i[5] ,
    \wbd_mbist8_dat_i[4] ,
    \wbd_mbist8_dat_i[3] ,
    \wbd_mbist8_dat_i[2] ,
    \wbd_mbist8_dat_i[1] ,
    \wbd_mbist8_dat_i[0] }),
    .wb_sel_i({\wbd_mbist8_sel_o[3] ,
    \wbd_mbist8_sel_o[2] ,
    \wbd_mbist8_sel_o[1] ,
    \wbd_mbist8_sel_o[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 u_sram1_2kb (.csb0(mem1_cen_b),
    .csb1(mem1_cen_a),
    .web0(mem1_web_b),
    .clk0(mem1_clk_b),
    .clk1(mem1_clk_a),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mem1_addr_b[10] ,
    \mem1_addr_b[9] ,
    \mem1_addr_b[8] ,
    \mem1_addr_b[7] ,
    \mem1_addr_b[6] ,
    \mem1_addr_b[5] ,
    \mem1_addr_b[4] ,
    \mem1_addr_b[3] ,
    \mem1_addr_b[2] }),
    .addr1({\mem1_addr_a[10] ,
    \mem1_addr_a[9] ,
    \mem1_addr_a[8] ,
    \mem1_addr_a[7] ,
    \mem1_addr_a[6] ,
    \mem1_addr_a[5] ,
    \mem1_addr_a[4] ,
    \mem1_addr_a[3] ,
    \mem1_addr_a[2] }),
    .din0({\mem1_din_b[31] ,
    \mem1_din_b[30] ,
    \mem1_din_b[29] ,
    \mem1_din_b[28] ,
    \mem1_din_b[27] ,
    \mem1_din_b[26] ,
    \mem1_din_b[25] ,
    \mem1_din_b[24] ,
    \mem1_din_b[23] ,
    \mem1_din_b[22] ,
    \mem1_din_b[21] ,
    \mem1_din_b[20] ,
    \mem1_din_b[19] ,
    \mem1_din_b[18] ,
    \mem1_din_b[17] ,
    \mem1_din_b[16] ,
    \mem1_din_b[15] ,
    \mem1_din_b[14] ,
    \mem1_din_b[13] ,
    \mem1_din_b[12] ,
    \mem1_din_b[11] ,
    \mem1_din_b[10] ,
    \mem1_din_b[9] ,
    \mem1_din_b[8] ,
    \mem1_din_b[7] ,
    \mem1_din_b[6] ,
    \mem1_din_b[5] ,
    \mem1_din_b[4] ,
    \mem1_din_b[3] ,
    \mem1_din_b[2] ,
    \mem1_din_b[1] ,
    \mem1_din_b[0] }),
    .dout0({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .dout1({\mem1_dout_a[31] ,
    \mem1_dout_a[30] ,
    \mem1_dout_a[29] ,
    \mem1_dout_a[28] ,
    \mem1_dout_a[27] ,
    \mem1_dout_a[26] ,
    \mem1_dout_a[25] ,
    \mem1_dout_a[24] ,
    \mem1_dout_a[23] ,
    \mem1_dout_a[22] ,
    \mem1_dout_a[21] ,
    \mem1_dout_a[20] ,
    \mem1_dout_a[19] ,
    \mem1_dout_a[18] ,
    \mem1_dout_a[17] ,
    \mem1_dout_a[16] ,
    \mem1_dout_a[15] ,
    \mem1_dout_a[14] ,
    \mem1_dout_a[13] ,
    \mem1_dout_a[12] ,
    \mem1_dout_a[11] ,
    \mem1_dout_a[10] ,
    \mem1_dout_a[9] ,
    \mem1_dout_a[8] ,
    \mem1_dout_a[7] ,
    \mem1_dout_a[6] ,
    \mem1_dout_a[5] ,
    \mem1_dout_a[4] ,
    \mem1_dout_a[3] ,
    \mem1_dout_a[2] ,
    \mem1_dout_a[1] ,
    \mem1_dout_a[0] }),
    .wmask0({\mem1_mask_b[3] ,
    \mem1_mask_b[2] ,
    \mem1_mask_b[1] ,
    \mem1_mask_b[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 u_sram2_2kb (.csb0(mem2_cen_b),
    .csb1(mem2_cen_a),
    .web0(mem2_web_b),
    .clk0(mem2_clk_b),
    .clk1(mem2_clk_a),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mem2_addr_b[10] ,
    \mem2_addr_b[9] ,
    \mem2_addr_b[8] ,
    \mem2_addr_b[7] ,
    \mem2_addr_b[6] ,
    \mem2_addr_b[5] ,
    \mem2_addr_b[4] ,
    \mem2_addr_b[3] ,
    \mem2_addr_b[2] }),
    .addr1({\mem2_addr_a[10] ,
    \mem2_addr_a[9] ,
    \mem2_addr_a[8] ,
    \mem2_addr_a[7] ,
    \mem2_addr_a[6] ,
    \mem2_addr_a[5] ,
    \mem2_addr_a[4] ,
    \mem2_addr_a[3] ,
    \mem2_addr_a[2] }),
    .din0({\mem2_din_b[31] ,
    \mem2_din_b[30] ,
    \mem2_din_b[29] ,
    \mem2_din_b[28] ,
    \mem2_din_b[27] ,
    \mem2_din_b[26] ,
    \mem2_din_b[25] ,
    \mem2_din_b[24] ,
    \mem2_din_b[23] ,
    \mem2_din_b[22] ,
    \mem2_din_b[21] ,
    \mem2_din_b[20] ,
    \mem2_din_b[19] ,
    \mem2_din_b[18] ,
    \mem2_din_b[17] ,
    \mem2_din_b[16] ,
    \mem2_din_b[15] ,
    \mem2_din_b[14] ,
    \mem2_din_b[13] ,
    \mem2_din_b[12] ,
    \mem2_din_b[11] ,
    \mem2_din_b[10] ,
    \mem2_din_b[9] ,
    \mem2_din_b[8] ,
    \mem2_din_b[7] ,
    \mem2_din_b[6] ,
    \mem2_din_b[5] ,
    \mem2_din_b[4] ,
    \mem2_din_b[3] ,
    \mem2_din_b[2] ,
    \mem2_din_b[1] ,
    \mem2_din_b[0] }),
    .dout0({_NC33,
    _NC34,
    _NC35,
    _NC36,
    _NC37,
    _NC38,
    _NC39,
    _NC40,
    _NC41,
    _NC42,
    _NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48,
    _NC49,
    _NC50,
    _NC51,
    _NC52,
    _NC53,
    _NC54,
    _NC55,
    _NC56,
    _NC57,
    _NC58,
    _NC59,
    _NC60,
    _NC61,
    _NC62,
    _NC63,
    _NC64}),
    .dout1({\mem2_dout_a[31] ,
    \mem2_dout_a[30] ,
    \mem2_dout_a[29] ,
    \mem2_dout_a[28] ,
    \mem2_dout_a[27] ,
    \mem2_dout_a[26] ,
    \mem2_dout_a[25] ,
    \mem2_dout_a[24] ,
    \mem2_dout_a[23] ,
    \mem2_dout_a[22] ,
    \mem2_dout_a[21] ,
    \mem2_dout_a[20] ,
    \mem2_dout_a[19] ,
    \mem2_dout_a[18] ,
    \mem2_dout_a[17] ,
    \mem2_dout_a[16] ,
    \mem2_dout_a[15] ,
    \mem2_dout_a[14] ,
    \mem2_dout_a[13] ,
    \mem2_dout_a[12] ,
    \mem2_dout_a[11] ,
    \mem2_dout_a[10] ,
    \mem2_dout_a[9] ,
    \mem2_dout_a[8] ,
    \mem2_dout_a[7] ,
    \mem2_dout_a[6] ,
    \mem2_dout_a[5] ,
    \mem2_dout_a[4] ,
    \mem2_dout_a[3] ,
    \mem2_dout_a[2] ,
    \mem2_dout_a[1] ,
    \mem2_dout_a[0] }),
    .wmask0({\mem2_mask_b[3] ,
    \mem2_mask_b[2] ,
    \mem2_mask_b[1] ,
    \mem2_mask_b[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 u_sram3_2kb (.csb0(mem3_cen_b),
    .csb1(mem3_cen_a),
    .web0(mem3_web_b),
    .clk0(mem3_clk_b),
    .clk1(mem3_clk_a),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mem3_addr_b[10] ,
    \mem3_addr_b[9] ,
    \mem3_addr_b[8] ,
    \mem3_addr_b[7] ,
    \mem3_addr_b[6] ,
    \mem3_addr_b[5] ,
    \mem3_addr_b[4] ,
    \mem3_addr_b[3] ,
    \mem3_addr_b[2] }),
    .addr1({\mem3_addr_a[10] ,
    \mem3_addr_a[9] ,
    \mem3_addr_a[8] ,
    \mem3_addr_a[7] ,
    \mem3_addr_a[6] ,
    \mem3_addr_a[5] ,
    \mem3_addr_a[4] ,
    \mem3_addr_a[3] ,
    \mem3_addr_a[2] }),
    .din0({\mem3_din_b[31] ,
    \mem3_din_b[30] ,
    \mem3_din_b[29] ,
    \mem3_din_b[28] ,
    \mem3_din_b[27] ,
    \mem3_din_b[26] ,
    \mem3_din_b[25] ,
    \mem3_din_b[24] ,
    \mem3_din_b[23] ,
    \mem3_din_b[22] ,
    \mem3_din_b[21] ,
    \mem3_din_b[20] ,
    \mem3_din_b[19] ,
    \mem3_din_b[18] ,
    \mem3_din_b[17] ,
    \mem3_din_b[16] ,
    \mem3_din_b[15] ,
    \mem3_din_b[14] ,
    \mem3_din_b[13] ,
    \mem3_din_b[12] ,
    \mem3_din_b[11] ,
    \mem3_din_b[10] ,
    \mem3_din_b[9] ,
    \mem3_din_b[8] ,
    \mem3_din_b[7] ,
    \mem3_din_b[6] ,
    \mem3_din_b[5] ,
    \mem3_din_b[4] ,
    \mem3_din_b[3] ,
    \mem3_din_b[2] ,
    \mem3_din_b[1] ,
    \mem3_din_b[0] }),
    .dout0({_NC65,
    _NC66,
    _NC67,
    _NC68,
    _NC69,
    _NC70,
    _NC71,
    _NC72,
    _NC73,
    _NC74,
    _NC75,
    _NC76,
    _NC77,
    _NC78,
    _NC79,
    _NC80,
    _NC81,
    _NC82,
    _NC83,
    _NC84,
    _NC85,
    _NC86,
    _NC87,
    _NC88,
    _NC89,
    _NC90,
    _NC91,
    _NC92,
    _NC93,
    _NC94,
    _NC95,
    _NC96}),
    .dout1({\mem3_dout_a[31] ,
    \mem3_dout_a[30] ,
    \mem3_dout_a[29] ,
    \mem3_dout_a[28] ,
    \mem3_dout_a[27] ,
    \mem3_dout_a[26] ,
    \mem3_dout_a[25] ,
    \mem3_dout_a[24] ,
    \mem3_dout_a[23] ,
    \mem3_dout_a[22] ,
    \mem3_dout_a[21] ,
    \mem3_dout_a[20] ,
    \mem3_dout_a[19] ,
    \mem3_dout_a[18] ,
    \mem3_dout_a[17] ,
    \mem3_dout_a[16] ,
    \mem3_dout_a[15] ,
    \mem3_dout_a[14] ,
    \mem3_dout_a[13] ,
    \mem3_dout_a[12] ,
    \mem3_dout_a[11] ,
    \mem3_dout_a[10] ,
    \mem3_dout_a[9] ,
    \mem3_dout_a[8] ,
    \mem3_dout_a[7] ,
    \mem3_dout_a[6] ,
    \mem3_dout_a[5] ,
    \mem3_dout_a[4] ,
    \mem3_dout_a[3] ,
    \mem3_dout_a[2] ,
    \mem3_dout_a[1] ,
    \mem3_dout_a[0] }),
    .wmask0({\mem3_mask_b[3] ,
    \mem3_mask_b[2] ,
    \mem3_mask_b[1] ,
    \mem3_mask_b[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 u_sram4_2kb (.csb0(mem4_cen_b),
    .csb1(mem4_cen_a),
    .web0(mem4_web_b),
    .clk0(mem4_clk_b),
    .clk1(mem4_clk_a),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mem4_addr_b[10] ,
    \mem4_addr_b[9] ,
    \mem4_addr_b[8] ,
    \mem4_addr_b[7] ,
    \mem4_addr_b[6] ,
    \mem4_addr_b[5] ,
    \mem4_addr_b[4] ,
    \mem4_addr_b[3] ,
    \mem4_addr_b[2] }),
    .addr1({\mem4_addr_a[10] ,
    \mem4_addr_a[9] ,
    \mem4_addr_a[8] ,
    \mem4_addr_a[7] ,
    \mem4_addr_a[6] ,
    \mem4_addr_a[5] ,
    \mem4_addr_a[4] ,
    \mem4_addr_a[3] ,
    \mem4_addr_a[2] }),
    .din0({\mem4_din_b[31] ,
    \mem4_din_b[30] ,
    \mem4_din_b[29] ,
    \mem4_din_b[28] ,
    \mem4_din_b[27] ,
    \mem4_din_b[26] ,
    \mem4_din_b[25] ,
    \mem4_din_b[24] ,
    \mem4_din_b[23] ,
    \mem4_din_b[22] ,
    \mem4_din_b[21] ,
    \mem4_din_b[20] ,
    \mem4_din_b[19] ,
    \mem4_din_b[18] ,
    \mem4_din_b[17] ,
    \mem4_din_b[16] ,
    \mem4_din_b[15] ,
    \mem4_din_b[14] ,
    \mem4_din_b[13] ,
    \mem4_din_b[12] ,
    \mem4_din_b[11] ,
    \mem4_din_b[10] ,
    \mem4_din_b[9] ,
    \mem4_din_b[8] ,
    \mem4_din_b[7] ,
    \mem4_din_b[6] ,
    \mem4_din_b[5] ,
    \mem4_din_b[4] ,
    \mem4_din_b[3] ,
    \mem4_din_b[2] ,
    \mem4_din_b[1] ,
    \mem4_din_b[0] }),
    .dout0({_NC97,
    _NC98,
    _NC99,
    _NC100,
    _NC101,
    _NC102,
    _NC103,
    _NC104,
    _NC105,
    _NC106,
    _NC107,
    _NC108,
    _NC109,
    _NC110,
    _NC111,
    _NC112,
    _NC113,
    _NC114,
    _NC115,
    _NC116,
    _NC117,
    _NC118,
    _NC119,
    _NC120,
    _NC121,
    _NC122,
    _NC123,
    _NC124,
    _NC125,
    _NC126,
    _NC127,
    _NC128}),
    .dout1({\mem4_dout_a[31] ,
    \mem4_dout_a[30] ,
    \mem4_dout_a[29] ,
    \mem4_dout_a[28] ,
    \mem4_dout_a[27] ,
    \mem4_dout_a[26] ,
    \mem4_dout_a[25] ,
    \mem4_dout_a[24] ,
    \mem4_dout_a[23] ,
    \mem4_dout_a[22] ,
    \mem4_dout_a[21] ,
    \mem4_dout_a[20] ,
    \mem4_dout_a[19] ,
    \mem4_dout_a[18] ,
    \mem4_dout_a[17] ,
    \mem4_dout_a[16] ,
    \mem4_dout_a[15] ,
    \mem4_dout_a[14] ,
    \mem4_dout_a[13] ,
    \mem4_dout_a[12] ,
    \mem4_dout_a[11] ,
    \mem4_dout_a[10] ,
    \mem4_dout_a[9] ,
    \mem4_dout_a[8] ,
    \mem4_dout_a[7] ,
    \mem4_dout_a[6] ,
    \mem4_dout_a[5] ,
    \mem4_dout_a[4] ,
    \mem4_dout_a[3] ,
    \mem4_dout_a[2] ,
    \mem4_dout_a[1] ,
    \mem4_dout_a[0] }),
    .wmask0({\mem4_mask_b[3] ,
    \mem4_mask_b[2] ,
    \mem4_mask_b[1] ,
    \mem4_mask_b[0] }));
 sky130_sram_1kbyte_1rw1r_32x256_8 u_sram5_1kb (.csb0(mem5_cen_b),
    .csb1(mem5_cen_a),
    .web0(mem5_web_b),
    .clk0(mem5_clk_b),
    .clk1(mem5_clk_a),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mem5_addr_b[9] ,
    \mem5_addr_b[8] ,
    \mem5_addr_b[7] ,
    \mem5_addr_b[6] ,
    \mem5_addr_b[5] ,
    \mem5_addr_b[4] ,
    \mem5_addr_b[3] ,
    \mem5_addr_b[2] }),
    .addr1({\mem5_addr_a[9] ,
    \mem5_addr_a[8] ,
    \mem5_addr_a[7] ,
    \mem5_addr_a[6] ,
    \mem5_addr_a[5] ,
    \mem5_addr_a[4] ,
    \mem5_addr_a[3] ,
    \mem5_addr_a[2] }),
    .din0({\mem5_din_b[31] ,
    \mem5_din_b[30] ,
    \mem5_din_b[29] ,
    \mem5_din_b[28] ,
    \mem5_din_b[27] ,
    \mem5_din_b[26] ,
    \mem5_din_b[25] ,
    \mem5_din_b[24] ,
    \mem5_din_b[23] ,
    \mem5_din_b[22] ,
    \mem5_din_b[21] ,
    \mem5_din_b[20] ,
    \mem5_din_b[19] ,
    \mem5_din_b[18] ,
    \mem5_din_b[17] ,
    \mem5_din_b[16] ,
    \mem5_din_b[15] ,
    \mem5_din_b[14] ,
    \mem5_din_b[13] ,
    \mem5_din_b[12] ,
    \mem5_din_b[11] ,
    \mem5_din_b[10] ,
    \mem5_din_b[9] ,
    \mem5_din_b[8] ,
    \mem5_din_b[7] ,
    \mem5_din_b[6] ,
    \mem5_din_b[5] ,
    \mem5_din_b[4] ,
    \mem5_din_b[3] ,
    \mem5_din_b[2] ,
    \mem5_din_b[1] ,
    \mem5_din_b[0] }),
    .dout0({_NC129,
    _NC130,
    _NC131,
    _NC132,
    _NC133,
    _NC134,
    _NC135,
    _NC136,
    _NC137,
    _NC138,
    _NC139,
    _NC140,
    _NC141,
    _NC142,
    _NC143,
    _NC144,
    _NC145,
    _NC146,
    _NC147,
    _NC148,
    _NC149,
    _NC150,
    _NC151,
    _NC152,
    _NC153,
    _NC154,
    _NC155,
    _NC156,
    _NC157,
    _NC158,
    _NC159,
    _NC160}),
    .dout1({\mem5_dout_a[31] ,
    \mem5_dout_a[30] ,
    \mem5_dout_a[29] ,
    \mem5_dout_a[28] ,
    \mem5_dout_a[27] ,
    \mem5_dout_a[26] ,
    \mem5_dout_a[25] ,
    \mem5_dout_a[24] ,
    \mem5_dout_a[23] ,
    \mem5_dout_a[22] ,
    \mem5_dout_a[21] ,
    \mem5_dout_a[20] ,
    \mem5_dout_a[19] ,
    \mem5_dout_a[18] ,
    \mem5_dout_a[17] ,
    \mem5_dout_a[16] ,
    \mem5_dout_a[15] ,
    \mem5_dout_a[14] ,
    \mem5_dout_a[13] ,
    \mem5_dout_a[12] ,
    \mem5_dout_a[11] ,
    \mem5_dout_a[10] ,
    \mem5_dout_a[9] ,
    \mem5_dout_a[8] ,
    \mem5_dout_a[7] ,
    \mem5_dout_a[6] ,
    \mem5_dout_a[5] ,
    \mem5_dout_a[4] ,
    \mem5_dout_a[3] ,
    \mem5_dout_a[2] ,
    \mem5_dout_a[1] ,
    \mem5_dout_a[0] }),
    .wmask0({\mem5_mask_b[3] ,
    \mem5_mask_b[2] ,
    \mem5_mask_b[1] ,
    \mem5_mask_b[0] }));
 sky130_sram_1kbyte_1rw1r_32x256_8 u_sram6_1kb (.csb0(mem6_cen_b),
    .csb1(mem6_cen_a),
    .web0(mem6_web_b),
    .clk0(mem6_clk_b),
    .clk1(mem6_clk_a),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mem6_addr_b[9] ,
    \mem6_addr_b[8] ,
    \mem6_addr_b[7] ,
    \mem6_addr_b[6] ,
    \mem6_addr_b[5] ,
    \mem6_addr_b[4] ,
    \mem6_addr_b[3] ,
    \mem6_addr_b[2] }),
    .addr1({\mem6_addr_a[9] ,
    \mem6_addr_a[8] ,
    \mem6_addr_a[7] ,
    \mem6_addr_a[6] ,
    \mem6_addr_a[5] ,
    \mem6_addr_a[4] ,
    \mem6_addr_a[3] ,
    \mem6_addr_a[2] }),
    .din0({\mem6_din_b[31] ,
    \mem6_din_b[30] ,
    \mem6_din_b[29] ,
    \mem6_din_b[28] ,
    \mem6_din_b[27] ,
    \mem6_din_b[26] ,
    \mem6_din_b[25] ,
    \mem6_din_b[24] ,
    \mem6_din_b[23] ,
    \mem6_din_b[22] ,
    \mem6_din_b[21] ,
    \mem6_din_b[20] ,
    \mem6_din_b[19] ,
    \mem6_din_b[18] ,
    \mem6_din_b[17] ,
    \mem6_din_b[16] ,
    \mem6_din_b[15] ,
    \mem6_din_b[14] ,
    \mem6_din_b[13] ,
    \mem6_din_b[12] ,
    \mem6_din_b[11] ,
    \mem6_din_b[10] ,
    \mem6_din_b[9] ,
    \mem6_din_b[8] ,
    \mem6_din_b[7] ,
    \mem6_din_b[6] ,
    \mem6_din_b[5] ,
    \mem6_din_b[4] ,
    \mem6_din_b[3] ,
    \mem6_din_b[2] ,
    \mem6_din_b[1] ,
    \mem6_din_b[0] }),
    .dout0({_NC161,
    _NC162,
    _NC163,
    _NC164,
    _NC165,
    _NC166,
    _NC167,
    _NC168,
    _NC169,
    _NC170,
    _NC171,
    _NC172,
    _NC173,
    _NC174,
    _NC175,
    _NC176,
    _NC177,
    _NC178,
    _NC179,
    _NC180,
    _NC181,
    _NC182,
    _NC183,
    _NC184,
    _NC185,
    _NC186,
    _NC187,
    _NC188,
    _NC189,
    _NC190,
    _NC191,
    _NC192}),
    .dout1({\mem6_dout_a[31] ,
    \mem6_dout_a[30] ,
    \mem6_dout_a[29] ,
    \mem6_dout_a[28] ,
    \mem6_dout_a[27] ,
    \mem6_dout_a[26] ,
    \mem6_dout_a[25] ,
    \mem6_dout_a[24] ,
    \mem6_dout_a[23] ,
    \mem6_dout_a[22] ,
    \mem6_dout_a[21] ,
    \mem6_dout_a[20] ,
    \mem6_dout_a[19] ,
    \mem6_dout_a[18] ,
    \mem6_dout_a[17] ,
    \mem6_dout_a[16] ,
    \mem6_dout_a[15] ,
    \mem6_dout_a[14] ,
    \mem6_dout_a[13] ,
    \mem6_dout_a[12] ,
    \mem6_dout_a[11] ,
    \mem6_dout_a[10] ,
    \mem6_dout_a[9] ,
    \mem6_dout_a[8] ,
    \mem6_dout_a[7] ,
    \mem6_dout_a[6] ,
    \mem6_dout_a[5] ,
    \mem6_dout_a[4] ,
    \mem6_dout_a[3] ,
    \mem6_dout_a[2] ,
    \mem6_dout_a[1] ,
    \mem6_dout_a[0] }),
    .wmask0({\mem6_mask_b[3] ,
    \mem6_mask_b[2] ,
    \mem6_mask_b[1] ,
    \mem6_mask_b[0] }));
 sky130_sram_1kbyte_1rw1r_32x256_8 u_sram7_1kb (.csb0(mem7_cen_b),
    .csb1(mem7_cen_a),
    .web0(mem7_web_b),
    .clk0(mem7_clk_b),
    .clk1(mem7_clk_a),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mem7_addr_b[9] ,
    \mem7_addr_b[8] ,
    \mem7_addr_b[7] ,
    \mem7_addr_b[6] ,
    \mem7_addr_b[5] ,
    \mem7_addr_b[4] ,
    \mem7_addr_b[3] ,
    \mem7_addr_b[2] }),
    .addr1({\mem7_addr_a[9] ,
    \mem7_addr_a[8] ,
    \mem7_addr_a[7] ,
    \mem7_addr_a[6] ,
    \mem7_addr_a[5] ,
    \mem7_addr_a[4] ,
    \mem7_addr_a[3] ,
    \mem7_addr_a[2] }),
    .din0({\mem7_din_b[31] ,
    \mem7_din_b[30] ,
    \mem7_din_b[29] ,
    \mem7_din_b[28] ,
    \mem7_din_b[27] ,
    \mem7_din_b[26] ,
    \mem7_din_b[25] ,
    \mem7_din_b[24] ,
    \mem7_din_b[23] ,
    \mem7_din_b[22] ,
    \mem7_din_b[21] ,
    \mem7_din_b[20] ,
    \mem7_din_b[19] ,
    \mem7_din_b[18] ,
    \mem7_din_b[17] ,
    \mem7_din_b[16] ,
    \mem7_din_b[15] ,
    \mem7_din_b[14] ,
    \mem7_din_b[13] ,
    \mem7_din_b[12] ,
    \mem7_din_b[11] ,
    \mem7_din_b[10] ,
    \mem7_din_b[9] ,
    \mem7_din_b[8] ,
    \mem7_din_b[7] ,
    \mem7_din_b[6] ,
    \mem7_din_b[5] ,
    \mem7_din_b[4] ,
    \mem7_din_b[3] ,
    \mem7_din_b[2] ,
    \mem7_din_b[1] ,
    \mem7_din_b[0] }),
    .dout0({_NC193,
    _NC194,
    _NC195,
    _NC196,
    _NC197,
    _NC198,
    _NC199,
    _NC200,
    _NC201,
    _NC202,
    _NC203,
    _NC204,
    _NC205,
    _NC206,
    _NC207,
    _NC208,
    _NC209,
    _NC210,
    _NC211,
    _NC212,
    _NC213,
    _NC214,
    _NC215,
    _NC216,
    _NC217,
    _NC218,
    _NC219,
    _NC220,
    _NC221,
    _NC222,
    _NC223,
    _NC224}),
    .dout1({\mem7_dout_a[31] ,
    \mem7_dout_a[30] ,
    \mem7_dout_a[29] ,
    \mem7_dout_a[28] ,
    \mem7_dout_a[27] ,
    \mem7_dout_a[26] ,
    \mem7_dout_a[25] ,
    \mem7_dout_a[24] ,
    \mem7_dout_a[23] ,
    \mem7_dout_a[22] ,
    \mem7_dout_a[21] ,
    \mem7_dout_a[20] ,
    \mem7_dout_a[19] ,
    \mem7_dout_a[18] ,
    \mem7_dout_a[17] ,
    \mem7_dout_a[16] ,
    \mem7_dout_a[15] ,
    \mem7_dout_a[14] ,
    \mem7_dout_a[13] ,
    \mem7_dout_a[12] ,
    \mem7_dout_a[11] ,
    \mem7_dout_a[10] ,
    \mem7_dout_a[9] ,
    \mem7_dout_a[8] ,
    \mem7_dout_a[7] ,
    \mem7_dout_a[6] ,
    \mem7_dout_a[5] ,
    \mem7_dout_a[4] ,
    \mem7_dout_a[3] ,
    \mem7_dout_a[2] ,
    \mem7_dout_a[1] ,
    \mem7_dout_a[0] }),
    .wmask0({\mem7_mask_b[3] ,
    \mem7_mask_b[2] ,
    \mem7_mask_b[1] ,
    \mem7_mask_b[0] }));
 sky130_sram_1kbyte_1rw1r_32x256_8 u_sram8_1kb (.csb0(mem8_cen_b),
    .csb1(mem8_cen_a),
    .web0(mem8_web_b),
    .clk0(mem8_clk_b),
    .clk1(mem8_clk_a),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mem8_addr_b[9] ,
    \mem8_addr_b[8] ,
    \mem8_addr_b[7] ,
    \mem8_addr_b[6] ,
    \mem8_addr_b[5] ,
    \mem8_addr_b[4] ,
    \mem8_addr_b[3] ,
    \mem8_addr_b[2] }),
    .addr1({\mem8_addr_a[9] ,
    \mem8_addr_a[8] ,
    \mem8_addr_a[7] ,
    \mem8_addr_a[6] ,
    \mem8_addr_a[5] ,
    \mem8_addr_a[4] ,
    \mem8_addr_a[3] ,
    \mem8_addr_a[2] }),
    .din0({\mem8_din_b[31] ,
    \mem8_din_b[30] ,
    \mem8_din_b[29] ,
    \mem8_din_b[28] ,
    \mem8_din_b[27] ,
    \mem8_din_b[26] ,
    \mem8_din_b[25] ,
    \mem8_din_b[24] ,
    \mem8_din_b[23] ,
    \mem8_din_b[22] ,
    \mem8_din_b[21] ,
    \mem8_din_b[20] ,
    \mem8_din_b[19] ,
    \mem8_din_b[18] ,
    \mem8_din_b[17] ,
    \mem8_din_b[16] ,
    \mem8_din_b[15] ,
    \mem8_din_b[14] ,
    \mem8_din_b[13] ,
    \mem8_din_b[12] ,
    \mem8_din_b[11] ,
    \mem8_din_b[10] ,
    \mem8_din_b[9] ,
    \mem8_din_b[8] ,
    \mem8_din_b[7] ,
    \mem8_din_b[6] ,
    \mem8_din_b[5] ,
    \mem8_din_b[4] ,
    \mem8_din_b[3] ,
    \mem8_din_b[2] ,
    \mem8_din_b[1] ,
    \mem8_din_b[0] }),
    .dout0({_NC225,
    _NC226,
    _NC227,
    _NC228,
    _NC229,
    _NC230,
    _NC231,
    _NC232,
    _NC233,
    _NC234,
    _NC235,
    _NC236,
    _NC237,
    _NC238,
    _NC239,
    _NC240,
    _NC241,
    _NC242,
    _NC243,
    _NC244,
    _NC245,
    _NC246,
    _NC247,
    _NC248,
    _NC249,
    _NC250,
    _NC251,
    _NC252,
    _NC253,
    _NC254,
    _NC255,
    _NC256}),
    .dout1({\mem8_dout_a[31] ,
    \mem8_dout_a[30] ,
    \mem8_dout_a[29] ,
    \mem8_dout_a[28] ,
    \mem8_dout_a[27] ,
    \mem8_dout_a[26] ,
    \mem8_dout_a[25] ,
    \mem8_dout_a[24] ,
    \mem8_dout_a[23] ,
    \mem8_dout_a[22] ,
    \mem8_dout_a[21] ,
    \mem8_dout_a[20] ,
    \mem8_dout_a[19] ,
    \mem8_dout_a[18] ,
    \mem8_dout_a[17] ,
    \mem8_dout_a[16] ,
    \mem8_dout_a[15] ,
    \mem8_dout_a[14] ,
    \mem8_dout_a[13] ,
    \mem8_dout_a[12] ,
    \mem8_dout_a[11] ,
    \mem8_dout_a[10] ,
    \mem8_dout_a[9] ,
    \mem8_dout_a[8] ,
    \mem8_dout_a[7] ,
    \mem8_dout_a[6] ,
    \mem8_dout_a[5] ,
    \mem8_dout_a[4] ,
    \mem8_dout_a[3] ,
    \mem8_dout_a[2] ,
    \mem8_dout_a[1] ,
    \mem8_dout_a[0] }),
    .wmask0({\mem8_mask_b[3] ,
    \mem8_mask_b[2] ,
    \mem8_mask_b[1] ,
    \mem8_mask_b[0] }));
 wb_host u_wb_host (.bist_rst_n(bist_rst_n),
    .lbist_clk_int(lbist_clk),
    .lbist_clk_out(lbist_clk),
    .scan_clk(scan_clk),
    .scan_en(scan_en),
    .scan_mode(scan_mode),
    .scan_rst_n(scan_rst_n),
    .user_clock1(wb_clk_i),
    .user_clock2(user_clock2),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbd_clk_int(wbd_clk_int),
    .wbd_clk_wh(wbd_clk_wh),
    .wbd_int_rst_n(wbd_int_rst_n),
    .wbm_ack_o(wbs_ack_o),
    .wbm_clk_i(wb_clk_i),
    .wbm_cyc_i(wbs_cyc_i),
    .wbm_rst_i(wb_rst_i),
    .wbm_stb_i(wbs_stb_i),
    .wbm_we_i(wbs_we_i),
    .wbs_ack_i(wbd_int_ack_o),
    .wbs_clk_i(wbd_clk_wh),
    .wbs_clk_out(wbd_clk_int),
    .wbs_cyc_o(wbd_int_cyc_i),
    .wbs_err_i(wbd_int_err_o),
    .wbs_stb_o(wbd_int_stb_i),
    .wbs_we_o(wbd_int_we_i),
    .cfg_clk_ctrl1({\cfg_clk_ctrl1[31] ,
    \cfg_clk_ctrl1[30] ,
    \cfg_clk_ctrl1[29] ,
    \cfg_clk_ctrl1[28] ,
    \cfg_clk_ctrl1[27] ,
    \cfg_clk_ctrl1[26] ,
    \cfg_clk_ctrl1[25] ,
    \cfg_clk_ctrl1[24] ,
    \cfg_clk_ctrl1[23] ,
    \cfg_clk_ctrl1[22] ,
    \cfg_clk_ctrl1[21] ,
    \cfg_clk_ctrl1[20] ,
    \cfg_clk_ctrl1[19] ,
    \cfg_clk_ctrl1[18] ,
    \cfg_clk_ctrl1[17] ,
    \cfg_clk_ctrl1[16] ,
    \cfg_clk_ctrl1[15] ,
    \cfg_clk_ctrl1[14] ,
    \cfg_clk_ctrl1[13] ,
    \cfg_clk_ctrl1[12] ,
    \cfg_clk_ctrl1[11] ,
    \cfg_clk_ctrl1[10] ,
    \cfg_clk_ctrl1[9] ,
    \cfg_clk_ctrl1[8] ,
    \cfg_clk_ctrl1[7] ,
    \cfg_clk_ctrl1[6] ,
    \cfg_clk_ctrl1[5] ,
    \cfg_clk_ctrl1[4] ,
    \cfg_clk_ctrl1[3] ,
    \cfg_clk_ctrl1[2] ,
    \cfg_clk_ctrl1[1] ,
    \cfg_clk_ctrl1[0] }),
    .cfg_clk_ctrl2({\cfg_clk_ctrl2[31] ,
    \cfg_clk_ctrl2[30] ,
    \cfg_clk_ctrl2[29] ,
    \cfg_clk_ctrl2[28] ,
    \cfg_clk_ctrl2[27] ,
    \cfg_clk_ctrl2[26] ,
    \cfg_clk_ctrl2[25] ,
    \cfg_clk_ctrl2[24] ,
    \cfg_clk_ctrl2[23] ,
    \cfg_clk_ctrl2[22] ,
    \cfg_clk_ctrl2[21] ,
    \cfg_clk_ctrl2[20] ,
    \cfg_clk_ctrl2[19] ,
    \cfg_clk_ctrl2[18] ,
    \cfg_clk_ctrl2[17] ,
    \cfg_clk_ctrl2[16] ,
    \cfg_clk_ctrl2[15] ,
    \cfg_clk_ctrl2[14] ,
    \cfg_clk_ctrl2[13] ,
    \cfg_clk_ctrl2[12] ,
    \cfg_clk_ctrl2[11] ,
    \cfg_clk_ctrl2[10] ,
    \cfg_clk_ctrl2[9] ,
    \cfg_clk_ctrl2[8] ,
    \cfg_clk_ctrl2[7] ,
    \cfg_clk_ctrl2[6] ,
    \cfg_clk_ctrl2[5] ,
    \cfg_clk_ctrl2[4] ,
    \cfg_clk_ctrl2[3] ,
    \cfg_clk_ctrl2[2] ,
    \cfg_clk_ctrl2[1] ,
    \cfg_clk_ctrl2[0] }),
    .cfg_cska_lbist({\cfg_clk_ctrl1[15] ,
    \cfg_clk_ctrl1[14] ,
    \cfg_clk_ctrl1[13] ,
    \cfg_clk_ctrl1[12] }),
    .cfg_cska_wh({\cfg_clk_ctrl1[3] ,
    \cfg_clk_ctrl1[2] ,
    \cfg_clk_ctrl1[1] ,
    \cfg_clk_ctrl1[0] }),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .la_data_out({la_data_out[127],
    la_data_out[126],
    la_data_out[125],
    la_data_out[124],
    la_data_out[123],
    la_data_out[122],
    la_data_out[121],
    la_data_out[120],
    la_data_out[119],
    la_data_out[118],
    la_data_out[117],
    la_data_out[116],
    la_data_out[115],
    la_data_out[114],
    la_data_out[113],
    la_data_out[112],
    la_data_out[111],
    la_data_out[110],
    la_data_out[109],
    la_data_out[108],
    la_data_out[107],
    la_data_out[106],
    la_data_out[105],
    la_data_out[104],
    la_data_out[103],
    la_data_out[102],
    la_data_out[101],
    la_data_out[100],
    la_data_out[99],
    la_data_out[98],
    la_data_out[97],
    la_data_out[96],
    la_data_out[95],
    la_data_out[94],
    la_data_out[93],
    la_data_out[92],
    la_data_out[91],
    la_data_out[90],
    la_data_out[89],
    la_data_out[88],
    la_data_out[87],
    la_data_out[86],
    la_data_out[85],
    la_data_out[84],
    la_data_out[83],
    la_data_out[82],
    la_data_out[81],
    la_data_out[80],
    la_data_out[79],
    la_data_out[78],
    la_data_out[77],
    la_data_out[76],
    la_data_out[75],
    la_data_out[74],
    la_data_out[73],
    la_data_out[72],
    la_data_out[71],
    la_data_out[70],
    la_data_out[69],
    la_data_out[68],
    la_data_out[67],
    la_data_out[66],
    la_data_out[65],
    la_data_out[64],
    la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32],
    la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}),
    .scan_in({\scan_in[7] ,
    \scan_in[6] ,
    \scan_in[5] ,
    \scan_in[4] ,
    \scan_in[3] ,
    \scan_in[2] ,
    \scan_in[1] ,
    \scan_in[0] }),
    .scan_out({\scan_out_mbist1[7] ,
    \scan_out_mbist1[6] ,
    \scan_out_mbist1[5] ,
    \scan_out_mbist1[4] ,
    \scan_out_mbist1[3] ,
    \scan_out_mbist1[2] ,
    \scan_out_mbist1[1] ,
    \scan_out_mbist1[0] }),
    .user_irq({user_irq[2],
    user_irq[1],
    user_irq[0]}),
    .wbm_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbm_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbm_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .wbm_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}),
    .wbs_adr_o({\wbd_int_adr_i[31] ,
    \wbd_int_adr_i[30] ,
    \wbd_int_adr_i[29] ,
    \wbd_int_adr_i[28] ,
    \wbd_int_adr_i[27] ,
    \wbd_int_adr_i[26] ,
    \wbd_int_adr_i[25] ,
    \wbd_int_adr_i[24] ,
    \wbd_int_adr_i[23] ,
    \wbd_int_adr_i[22] ,
    \wbd_int_adr_i[21] ,
    \wbd_int_adr_i[20] ,
    \wbd_int_adr_i[19] ,
    \wbd_int_adr_i[18] ,
    \wbd_int_adr_i[17] ,
    \wbd_int_adr_i[16] ,
    \wbd_int_adr_i[15] ,
    \wbd_int_adr_i[14] ,
    \wbd_int_adr_i[13] ,
    \wbd_int_adr_i[12] ,
    \wbd_int_adr_i[11] ,
    \wbd_int_adr_i[10] ,
    \wbd_int_adr_i[9] ,
    \wbd_int_adr_i[8] ,
    \wbd_int_adr_i[7] ,
    \wbd_int_adr_i[6] ,
    \wbd_int_adr_i[5] ,
    \wbd_int_adr_i[4] ,
    \wbd_int_adr_i[3] ,
    \wbd_int_adr_i[2] ,
    \wbd_int_adr_i[1] ,
    \wbd_int_adr_i[0] }),
    .wbs_dat_i({\wbd_int_dat_o[31] ,
    \wbd_int_dat_o[30] ,
    \wbd_int_dat_o[29] ,
    \wbd_int_dat_o[28] ,
    \wbd_int_dat_o[27] ,
    \wbd_int_dat_o[26] ,
    \wbd_int_dat_o[25] ,
    \wbd_int_dat_o[24] ,
    \wbd_int_dat_o[23] ,
    \wbd_int_dat_o[22] ,
    \wbd_int_dat_o[21] ,
    \wbd_int_dat_o[20] ,
    \wbd_int_dat_o[19] ,
    \wbd_int_dat_o[18] ,
    \wbd_int_dat_o[17] ,
    \wbd_int_dat_o[16] ,
    \wbd_int_dat_o[15] ,
    \wbd_int_dat_o[14] ,
    \wbd_int_dat_o[13] ,
    \wbd_int_dat_o[12] ,
    \wbd_int_dat_o[11] ,
    \wbd_int_dat_o[10] ,
    \wbd_int_dat_o[9] ,
    \wbd_int_dat_o[8] ,
    \wbd_int_dat_o[7] ,
    \wbd_int_dat_o[6] ,
    \wbd_int_dat_o[5] ,
    \wbd_int_dat_o[4] ,
    \wbd_int_dat_o[3] ,
    \wbd_int_dat_o[2] ,
    \wbd_int_dat_o[1] ,
    \wbd_int_dat_o[0] }),
    .wbs_dat_o({\wbd_int_dat_i[31] ,
    \wbd_int_dat_i[30] ,
    \wbd_int_dat_i[29] ,
    \wbd_int_dat_i[28] ,
    \wbd_int_dat_i[27] ,
    \wbd_int_dat_i[26] ,
    \wbd_int_dat_i[25] ,
    \wbd_int_dat_i[24] ,
    \wbd_int_dat_i[23] ,
    \wbd_int_dat_i[22] ,
    \wbd_int_dat_i[21] ,
    \wbd_int_dat_i[20] ,
    \wbd_int_dat_i[19] ,
    \wbd_int_dat_i[18] ,
    \wbd_int_dat_i[17] ,
    \wbd_int_dat_i[16] ,
    \wbd_int_dat_i[15] ,
    \wbd_int_dat_i[14] ,
    \wbd_int_dat_i[13] ,
    \wbd_int_dat_i[12] ,
    \wbd_int_dat_i[11] ,
    \wbd_int_dat_i[10] ,
    \wbd_int_dat_i[9] ,
    \wbd_int_dat_i[8] ,
    \wbd_int_dat_i[7] ,
    \wbd_int_dat_i[6] ,
    \wbd_int_dat_i[5] ,
    \wbd_int_dat_i[4] ,
    \wbd_int_dat_i[3] ,
    \wbd_int_dat_i[2] ,
    \wbd_int_dat_i[1] ,
    \wbd_int_dat_i[0] }),
    .wbs_sel_o({\wbd_int_sel_i[3] ,
    \wbd_int_sel_i[2] ,
    \wbd_int_sel_i[1] ,
    \wbd_int_sel_i[0] }));
endmodule
