///////////////////////////////////////////////////////////////////////
// SPDX-FileCopyrightText: 2021 , Dinesh Annayya                          
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0
// SPDX-FileContributor: Created by Dinesh Annayya <dinesha@opencores.org>
//
//////////////////////////////////////////////////////////////////////
//------------------------------------------------------------------------
// This module is used to generate 1us based on config value
//------------------------------------------------------------------------

module pulse_gen_type2 #(parameter WD = 10)
    (
	output logic           clk_pulse,

	input logic            clk,
        input logic            reset_n,
	input logic [WD-1:0]   cfg_max_cnt
);


logic [WD-1:0]  cnt;


always @ (posedge clk or negedge reset_n)
begin
   if (reset_n == 1'b0) begin 
      cnt <= 'b0;
      clk_pulse <= 'b0;
   end else begin 
      if(cnt == cfg_max_cnt) begin
          cnt       <= 0;
          clk_pulse <= 1'b1;
      end else begin
          cnt       <= cnt +1;
          clk_pulse <= 1'b0;
      end
   end
end

endmodule

